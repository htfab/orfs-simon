module ttsimon (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire net26;
 wire net25;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire net24;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire net23;
 wire net22;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire net21;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire net20;
 wire _0312_;
 wire net19;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire net18;
 wire net17;
 wire net16;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire net15;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire net14;
 wire _0436_;
 wire _0437_;
 wire net13;
 wire _0439_;
 wire _0440_;
 wire net12;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire net11;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire net10;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire net9;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire net8;
 wire net7;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire net6;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire net5;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire net4;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire net3;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire net2;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire net135;
 wire net134;
 wire net133;
 wire _0749_;
 wire net132;
 wire _0751_;
 wire _0752_;
 wire net131;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire net130;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire net129;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire net128;
 wire net127;
 wire net126;
 wire net125;
 wire _0793_;
 wire _0794_;
 wire net124;
 wire _0796_;
 wire net123;
 wire net122;
 wire net121;
 wire net120;
 wire net119;
 wire net118;
 wire net117;
 wire net116;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire net115;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire net114;
 wire _0818_;
 wire net113;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire net112;
 wire _0832_;
 wire _0833_;
 wire net111;
 wire _0835_;
 wire net110;
 wire net109;
 wire net108;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire net107;
 wire _0845_;
 wire net106;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire net105;
 wire net104;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire net103;
 wire net102;
 wire _0862_;
 wire net100;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire net99;
 wire _0871_;
 wire net98;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire net93;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire net92;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire net91;
 wire _0910_;
 wire net90;
 wire _0912_;
 wire net89;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire net88;
 wire net87;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire net86;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire net85;
 wire _0940_;
 wire _0941_;
 wire net84;
 wire net83;
 wire _0944_;
 wire _0945_;
 wire net82;
 wire net81;
 wire _0948_;
 wire _0949_;
 wire net80;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire net79;
 wire net78;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire net77;
 wire net76;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire net75;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire net74;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire net73;
 wire net72;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire net71;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire net70;
 wire _1008_;
 wire _1009_;
 wire net69;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire net68;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire net67;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire net66;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire net65;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire net64;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire net63;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire net62;
 wire _1102_;
 wire net61;
 wire net60;
 wire net59;
 wire _1106_;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire _1111_;
 wire _1112_;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire net50;
 wire _1121_;
 wire net49;
 wire net48;
 wire _1124_;
 wire net47;
 wire net46;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire net45;
 wire net44;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire net43;
 wire _1136_;
 wire net42;
 wire net41;
 wire _1139_;
 wire net40;
 wire net39;
 wire _1142_;
 wire net38;
 wire net37;
 wire _1145_;
 wire net36;
 wire net35;
 wire net34;
 wire _1149_;
 wire _1150_;
 wire net33;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire net32;
 wire _1161_;
 wire net31;
 wire net30;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire net29;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire net28;
 wire _1210_;
 wire net27;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire net1;
 wire \simon1.millis_counter[0] ;
 wire \simon1.millis_counter[1] ;
 wire \simon1.millis_counter[2] ;
 wire \simon1.millis_counter[3] ;
 wire \simon1.millis_counter[4] ;
 wire \simon1.millis_counter[5] ;
 wire \simon1.millis_counter[6] ;
 wire \simon1.millis_counter[7] ;
 wire \simon1.millis_counter[8] ;
 wire \simon1.millis_counter[9] ;
 wire \simon1.next_random[0] ;
 wire \simon1.next_random[1] ;
 wire \simon1.play1.freq[0] ;
 wire \simon1.play1.freq[1] ;
 wire \simon1.play1.freq[2] ;
 wire \simon1.play1.freq[3] ;
 wire \simon1.play1.freq[4] ;
 wire \simon1.play1.freq[5] ;
 wire \simon1.play1.freq[6] ;
 wire \simon1.play1.freq[7] ;
 wire \simon1.play1.freq[8] ;
 wire \simon1.play1.freq[9] ;
 wire \simon1.play1.tick_counter[0] ;
 wire \simon1.play1.tick_counter[10] ;
 wire \simon1.play1.tick_counter[11] ;
 wire \simon1.play1.tick_counter[12] ;
 wire \simon1.play1.tick_counter[13] ;
 wire \simon1.play1.tick_counter[14] ;
 wire \simon1.play1.tick_counter[15] ;
 wire \simon1.play1.tick_counter[16] ;
 wire \simon1.play1.tick_counter[17] ;
 wire \simon1.play1.tick_counter[18] ;
 wire \simon1.play1.tick_counter[19] ;
 wire \simon1.play1.tick_counter[1] ;
 wire \simon1.play1.tick_counter[20] ;
 wire \simon1.play1.tick_counter[21] ;
 wire \simon1.play1.tick_counter[22] ;
 wire \simon1.play1.tick_counter[23] ;
 wire \simon1.play1.tick_counter[24] ;
 wire \simon1.play1.tick_counter[25] ;
 wire \simon1.play1.tick_counter[26] ;
 wire \simon1.play1.tick_counter[27] ;
 wire \simon1.play1.tick_counter[28] ;
 wire \simon1.play1.tick_counter[29] ;
 wire \simon1.play1.tick_counter[2] ;
 wire \simon1.play1.tick_counter[30] ;
 wire \simon1.play1.tick_counter[31] ;
 wire \simon1.play1.tick_counter[3] ;
 wire \simon1.play1.tick_counter[4] ;
 wire \simon1.play1.tick_counter[5] ;
 wire \simon1.play1.tick_counter[6] ;
 wire \simon1.play1.tick_counter[7] ;
 wire \simon1.play1.tick_counter[8] ;
 wire \simon1.play1.tick_counter[9] ;
 wire \simon1.score1.active_digit ;
 wire \simon1.score1.ena ;
 wire \simon1.score1.inc ;
 wire \simon1.score1.ones[0] ;
 wire \simon1.score1.ones[1] ;
 wire \simon1.score1.ones[2] ;
 wire \simon1.score1.ones[3] ;
 wire \simon1.score1.tens[0] ;
 wire \simon1.score1.tens[1] ;
 wire \simon1.score1.tens[2] ;
 wire \simon1.score1.tens[3] ;
 wire \simon1.score_rst ;
 wire \simon1.seq[0][0] ;
 wire \simon1.seq[0][1] ;
 wire \simon1.seq[10][0] ;
 wire \simon1.seq[10][1] ;
 wire \simon1.seq[11][0] ;
 wire \simon1.seq[11][1] ;
 wire \simon1.seq[12][0] ;
 wire \simon1.seq[12][1] ;
 wire \simon1.seq[13][0] ;
 wire \simon1.seq[13][1] ;
 wire \simon1.seq[14][0] ;
 wire \simon1.seq[14][1] ;
 wire \simon1.seq[15][0] ;
 wire \simon1.seq[15][1] ;
 wire \simon1.seq[16][0] ;
 wire \simon1.seq[16][1] ;
 wire \simon1.seq[17][0] ;
 wire \simon1.seq[17][1] ;
 wire \simon1.seq[18][0] ;
 wire \simon1.seq[18][1] ;
 wire \simon1.seq[19][0] ;
 wire \simon1.seq[19][1] ;
 wire \simon1.seq[1][0] ;
 wire \simon1.seq[1][1] ;
 wire \simon1.seq[20][0] ;
 wire \simon1.seq[20][1] ;
 wire \simon1.seq[21][0] ;
 wire \simon1.seq[21][1] ;
 wire \simon1.seq[22][0] ;
 wire \simon1.seq[22][1] ;
 wire \simon1.seq[23][0] ;
 wire \simon1.seq[23][1] ;
 wire \simon1.seq[24][0] ;
 wire \simon1.seq[24][1] ;
 wire \simon1.seq[25][0] ;
 wire \simon1.seq[25][1] ;
 wire \simon1.seq[26][0] ;
 wire \simon1.seq[26][1] ;
 wire \simon1.seq[27][0] ;
 wire \simon1.seq[27][1] ;
 wire \simon1.seq[28][0] ;
 wire \simon1.seq[28][1] ;
 wire \simon1.seq[29][0] ;
 wire \simon1.seq[29][1] ;
 wire \simon1.seq[2][0] ;
 wire \simon1.seq[2][1] ;
 wire \simon1.seq[30][0] ;
 wire \simon1.seq[30][1] ;
 wire \simon1.seq[31][0] ;
 wire \simon1.seq[31][1] ;
 wire \simon1.seq[3][0] ;
 wire \simon1.seq[3][1] ;
 wire \simon1.seq[4][0] ;
 wire \simon1.seq[4][1] ;
 wire \simon1.seq[5][0] ;
 wire \simon1.seq[5][1] ;
 wire \simon1.seq[6][0] ;
 wire \simon1.seq[6][1] ;
 wire \simon1.seq[7][0] ;
 wire \simon1.seq[7][1] ;
 wire \simon1.seq[8][0] ;
 wire \simon1.seq[8][1] ;
 wire \simon1.seq[9][0] ;
 wire \simon1.seq[9][1] ;
 wire \simon1.seq_counter[0] ;
 wire \simon1.seq_counter[1] ;
 wire \simon1.seq_counter[2] ;
 wire \simon1.seq_counter[3] ;
 wire \simon1.seq_counter[4] ;
 wire \simon1.seq_length[0] ;
 wire \simon1.seq_length[1] ;
 wire \simon1.seq_length[2] ;
 wire \simon1.seq_length[3] ;
 wire \simon1.seq_length[4] ;
 wire \simon1.state[0] ;
 wire \simon1.state[1] ;
 wire \simon1.state[2] ;
 wire \simon1.state[3] ;
 wire \simon1.state[4] ;
 wire \simon1.state[5] ;
 wire \simon1.state[6] ;
 wire \simon1.state[7] ;
 wire \simon1.tick_counter[0] ;
 wire \simon1.tick_counter[10] ;
 wire \simon1.tick_counter[11] ;
 wire \simon1.tick_counter[12] ;
 wire \simon1.tick_counter[13] ;
 wire \simon1.tick_counter[14] ;
 wire \simon1.tick_counter[15] ;
 wire \simon1.tick_counter[1] ;
 wire \simon1.tick_counter[2] ;
 wire \simon1.tick_counter[3] ;
 wire \simon1.tick_counter[4] ;
 wire \simon1.tick_counter[5] ;
 wire \simon1.tick_counter[6] ;
 wire \simon1.tick_counter[7] ;
 wire \simon1.tick_counter[8] ;
 wire \simon1.tick_counter[9] ;
 wire \simon1.tone_sequence_counter[0] ;
 wire \simon1.tone_sequence_counter[1] ;
 wire \simon1.tone_sequence_counter[2] ;
 wire \simon1.user_input[0] ;
 wire \simon1.user_input[1] ;
 wire clknet_0_clk;
 wire net101;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_tiehi \simon1.play1.tick_counter[10]$_SDFFE_PN0N__137  (.L_HI(net137));
 sg13g2_tiehi \simon1.play1.tick_counter[0]$_SDFFE_PN0N__136  (.L_HI(net136));
 sg13g2_tiehi \simon1.play1.sound$_SDFFE_PP0N__135  (.L_HI(net135));
 sg13g2_nand2b_1 _1403_ (.Y(_0749_),
    .B(\simon1.score1.ones[1] ),
    .A_N(net71));
 sg13g2_tiehi \simon1.play1.freq[9]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_nand2_1 _1405_ (.Y(_0751_),
    .A(net71),
    .B(\simon1.score1.tens[1] ));
 sg13g2_nand3_1 _1406_ (.B(_0749_),
    .C(_0751_),
    .A(\simon1.score1.ena ),
    .Y(_0752_));
 sg13g2_tiehi \simon1.play1.freq[8]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_inv_1 _1408_ (.Y(_0754_),
    .A(_0752_));
 sg13g2_inv_1 _1409_ (.Y(_0755_),
    .A(\simon1.score1.tens[2] ));
 sg13g2_nor2_1 _1410_ (.A(net71),
    .B(\simon1.score1.ones[2] ),
    .Y(_0756_));
 sg13g2_a21oi_1 _1411_ (.A1(net71),
    .A2(_0755_),
    .Y(_0757_),
    .B1(_0756_));
 sg13g2_or2_2 _1412_ (.X(_0758_),
    .B(_0757_),
    .A(_0026_));
 sg13g2_tiehi \simon1.play1.freq[7]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_inv_1 _1414_ (.Y(_0760_),
    .A(\simon1.score1.ones[3] ));
 sg13g2_nand2_1 _1415_ (.Y(_0761_),
    .A(net71),
    .B(\simon1.score1.tens[3] ));
 sg13g2_o21ai_1 _1416_ (.B1(_0761_),
    .Y(_0762_),
    .A1(net71),
    .A2(_0760_));
 sg13g2_nor3_1 _1417_ (.A(_0026_),
    .B(_0762_),
    .C(_0757_),
    .Y(_0763_));
 sg13g2_nand2b_1 _1418_ (.Y(_0764_),
    .B(\simon1.score1.ones[0] ),
    .A_N(net71));
 sg13g2_nand2_1 _1419_ (.Y(_0765_),
    .A(\simon1.score1.tens[0] ),
    .B(net71));
 sg13g2_nand3_1 _1420_ (.B(_0764_),
    .C(_0765_),
    .A(\simon1.score1.ena ),
    .Y(_0766_));
 sg13g2_tiehi \simon1.play1.freq[6]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_mux2_1 _1422_ (.A0(_0758_),
    .A1(_0763_),
    .S(_0766_),
    .X(_0768_));
 sg13g2_nor2_2 _1423_ (.A(_0026_),
    .B(_0762_),
    .Y(_0769_));
 sg13g2_nor2_2 _1424_ (.A(_0758_),
    .B(_0752_),
    .Y(_0770_));
 sg13g2_nor2_1 _1425_ (.A(_0769_),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_a21oi_1 _1426_ (.A1(_0754_),
    .A2(_0768_),
    .Y(_0772_),
    .B1(_0771_));
 sg13g2_xor2_1 _1427_ (.B(_0772_),
    .A(net6),
    .X(_0204_));
 sg13g2_xor2_1 _1428_ (.B(_0766_),
    .A(_0752_),
    .X(_0773_));
 sg13g2_a21oi_1 _1429_ (.A1(_0758_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0771_));
 sg13g2_xor2_1 _1430_ (.B(_0774_),
    .A(net6),
    .X(_0205_));
 sg13g2_o21ai_1 _1431_ (.B1(_0769_),
    .Y(_0775_),
    .A1(_0758_),
    .A2(_0766_));
 sg13g2_nor2b_1 _1432_ (.A(_0770_),
    .B_N(_0775_),
    .Y(_0776_));
 sg13g2_xnor2_1 _1433_ (.Y(_0206_),
    .A(net6),
    .B(_0776_));
 sg13g2_nand2_1 _1434_ (.Y(_0777_),
    .A(_0758_),
    .B(_0752_));
 sg13g2_nand2_1 _1435_ (.Y(_0778_),
    .A(_0769_),
    .B(_0770_));
 sg13g2_nand2_1 _1436_ (.Y(_0779_),
    .A(_0777_),
    .B(_0778_));
 sg13g2_nor2_1 _1437_ (.A(_0752_),
    .B(_0766_),
    .Y(_0780_));
 sg13g2_a221oi_1 _1438_ (.B2(_0758_),
    .C1(_0771_),
    .B1(_0780_),
    .A1(_0766_),
    .Y(_0781_),
    .A2(_0779_));
 sg13g2_xor2_1 _1439_ (.B(_0781_),
    .A(net6),
    .X(_0207_));
 sg13g2_a21oi_1 _1440_ (.A1(_0769_),
    .A2(_0752_),
    .Y(_0782_),
    .B1(_0770_));
 sg13g2_nor2_1 _1441_ (.A(_0766_),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_xor2_1 _1442_ (.B(_0783_),
    .A(net6),
    .X(_0208_));
 sg13g2_and2_1 _1443_ (.A(_0769_),
    .B(_0758_),
    .X(_0784_));
 sg13g2_o21ai_1 _1444_ (.B1(_0766_),
    .Y(_0785_),
    .A1(_0752_),
    .A2(_0763_));
 sg13g2_o21ai_1 _1445_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0770_),
    .A2(_0784_));
 sg13g2_xnor2_1 _1446_ (.Y(_0209_),
    .A(net6),
    .B(_0786_));
 sg13g2_nand3_1 _1447_ (.B(_0752_),
    .C(_0766_),
    .A(_0758_),
    .Y(_0787_));
 sg13g2_nand3b_1 _1448_ (.B(_0778_),
    .C(_0787_),
    .Y(_0788_),
    .A_N(_0771_));
 sg13g2_xnor2_1 _1449_ (.Y(_0210_),
    .A(net6),
    .B(_0788_));
 sg13g2_tiehi \simon1.play1.freq[5]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \simon1.play1.freq[4]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \simon1.play1.freq[3]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \simon1.play1.freq[2]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_nor3_2 _1454_ (.A(net3),
    .B(net4),
    .C(net5),
    .Y(_0793_));
 sg13g2_nor2b_2 _1455_ (.A(net2),
    .B_N(_0793_),
    .Y(_0794_));
 sg13g2_tiehi \simon1.play1.freq[1]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_inv_1 _1457_ (.Y(_0796_),
    .A(net96));
 sg13g2_tiehi \simon1.play1.freq[0]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \simon1.next_random[1]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_a21o_1 _1460_ (.A2(_0794_),
    .A1(\simon1.state[0] ),
    .B1(net94),
    .X(_0005_));
 sg13g2_tiehi \simon1.next_random[0]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \simon1.millis_counter[9]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \simon1.millis_counter[8]$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \simon1.millis_counter[7]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \simon1.millis_counter[6]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \simon1.millis_counter[5]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_mux4_1 _1467_ (.S0(net85),
    .A0(\simon1.seq[0][0] ),
    .A1(\simon1.seq[1][0] ),
    .A2(\simon1.seq[2][0] ),
    .A3(\simon1.seq[3][0] ),
    .S1(net83),
    .X(_0805_));
 sg13g2_mux4_1 _1468_ (.S0(net85),
    .A0(\simon1.seq[4][0] ),
    .A1(\simon1.seq[5][0] ),
    .A2(\simon1.seq[6][0] ),
    .A3(\simon1.seq[7][0] ),
    .S1(net83),
    .X(_0806_));
 sg13g2_mux4_1 _1469_ (.S0(net85),
    .A0(\simon1.seq[8][0] ),
    .A1(\simon1.seq[9][0] ),
    .A2(\simon1.seq[10][0] ),
    .A3(\simon1.seq[11][0] ),
    .S1(net83),
    .X(_0807_));
 sg13g2_mux4_1 _1470_ (.S0(net85),
    .A0(\simon1.seq[12][0] ),
    .A1(\simon1.seq[13][0] ),
    .A2(\simon1.seq[14][0] ),
    .A3(\simon1.seq[15][0] ),
    .S1(net83),
    .X(_0808_));
 sg13g2_tiehi \simon1.millis_counter[4]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_mux4_1 _1472_ (.S0(_0002_),
    .A0(_0805_),
    .A1(_0806_),
    .A2(_0807_),
    .A3(_0808_),
    .S1(_0003_),
    .X(_0810_));
 sg13g2_mux4_1 _1473_ (.S0(net84),
    .A0(\simon1.seq[16][0] ),
    .A1(\simon1.seq[17][0] ),
    .A2(\simon1.seq[18][0] ),
    .A3(\simon1.seq[19][0] ),
    .S1(net82),
    .X(_0811_));
 sg13g2_mux4_1 _1474_ (.S0(net84),
    .A0(\simon1.seq[20][0] ),
    .A1(\simon1.seq[21][0] ),
    .A2(\simon1.seq[22][0] ),
    .A3(\simon1.seq[23][0] ),
    .S1(net82),
    .X(_0812_));
 sg13g2_mux4_1 _1475_ (.S0(net84),
    .A0(\simon1.seq[24][0] ),
    .A1(\simon1.seq[25][0] ),
    .A2(\simon1.seq[26][0] ),
    .A3(\simon1.seq[27][0] ),
    .S1(net82),
    .X(_0813_));
 sg13g2_mux4_1 _1476_ (.S0(net84),
    .A0(\simon1.seq[28][0] ),
    .A1(\simon1.seq[29][0] ),
    .A2(\simon1.seq[30][0] ),
    .A3(\simon1.seq[31][0] ),
    .S1(net82),
    .X(_0814_));
 sg13g2_mux4_1 _1477_ (.S0(_0002_),
    .A0(_0811_),
    .A1(_0812_),
    .A2(_0813_),
    .A3(_0814_),
    .S1(_0003_),
    .X(_0815_));
 sg13g2_mux2_1 _1478_ (.A0(_0810_),
    .A1(_0815_),
    .S(_0004_),
    .X(_0816_));
 sg13g2_tiehi \simon1.millis_counter[3]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_xnor2_1 _1480_ (.Y(_0818_),
    .A(\simon1.user_input[0] ),
    .B(net44));
 sg13g2_tiehi \simon1.millis_counter[2]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_mux4_1 _1482_ (.S0(net85),
    .A0(\simon1.seq[0][1] ),
    .A1(\simon1.seq[1][1] ),
    .A2(\simon1.seq[2][1] ),
    .A3(\simon1.seq[3][1] ),
    .S1(net83),
    .X(_0820_));
 sg13g2_mux4_1 _1483_ (.S0(net85),
    .A0(\simon1.seq[4][1] ),
    .A1(\simon1.seq[5][1] ),
    .A2(\simon1.seq[6][1] ),
    .A3(\simon1.seq[7][1] ),
    .S1(net83),
    .X(_0821_));
 sg13g2_mux4_1 _1484_ (.S0(net85),
    .A0(\simon1.seq[8][1] ),
    .A1(\simon1.seq[9][1] ),
    .A2(\simon1.seq[10][1] ),
    .A3(\simon1.seq[11][1] ),
    .S1(net83),
    .X(_0822_));
 sg13g2_mux4_1 _1485_ (.S0(net85),
    .A0(\simon1.seq[12][1] ),
    .A1(\simon1.seq[13][1] ),
    .A2(\simon1.seq[14][1] ),
    .A3(\simon1.seq[15][1] ),
    .S1(net83),
    .X(_0823_));
 sg13g2_mux4_1 _1486_ (.S0(_0002_),
    .A0(_0820_),
    .A1(_0821_),
    .A2(_0822_),
    .A3(_0823_),
    .S1(_0003_),
    .X(_0824_));
 sg13g2_mux4_1 _1487_ (.S0(net84),
    .A0(\simon1.seq[16][1] ),
    .A1(\simon1.seq[17][1] ),
    .A2(\simon1.seq[18][1] ),
    .A3(\simon1.seq[19][1] ),
    .S1(net82),
    .X(_0825_));
 sg13g2_mux4_1 _1488_ (.S0(net84),
    .A0(\simon1.seq[20][1] ),
    .A1(\simon1.seq[21][1] ),
    .A2(\simon1.seq[22][1] ),
    .A3(\simon1.seq[23][1] ),
    .S1(net82),
    .X(_0826_));
 sg13g2_mux4_1 _1489_ (.S0(net84),
    .A0(\simon1.seq[24][1] ),
    .A1(\simon1.seq[25][1] ),
    .A2(\simon1.seq[26][1] ),
    .A3(\simon1.seq[27][1] ),
    .S1(net82),
    .X(_0827_));
 sg13g2_mux4_1 _1490_ (.S0(net84),
    .A0(\simon1.seq[28][1] ),
    .A1(\simon1.seq[29][1] ),
    .A2(\simon1.seq[30][1] ),
    .A3(\simon1.seq[31][1] ),
    .S1(net82),
    .X(_0828_));
 sg13g2_mux4_1 _1491_ (.S0(_0002_),
    .A0(_0825_),
    .A1(_0826_),
    .A2(_0827_),
    .A3(_0828_),
    .S1(_0003_),
    .X(_0829_));
 sg13g2_mux2_2 _1492_ (.A0(_0824_),
    .A1(_0829_),
    .S(_0004_),
    .X(_0830_));
 sg13g2_tiehi \simon1.millis_counter[1]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_xnor2_1 _1494_ (.Y(_0832_),
    .A(\simon1.user_input[1] ),
    .B(_0830_));
 sg13g2_nand2_2 _1495_ (.Y(_0833_),
    .A(_0818_),
    .B(_0832_));
 sg13g2_tiehi \simon1.millis_counter[0]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_inv_2 _1497_ (.Y(_0835_),
    .A(net61));
 sg13g2_tiehi _2618__112 (.L_HI(net112));
 sg13g2_tiehi _2617__111 (.L_HI(net111));
 sg13g2_tiehi _2616__110 (.L_HI(net110));
 sg13g2_nand2b_1 _1501_ (.Y(_0839_),
    .B(\simon1.millis_counter[8] ),
    .A_N(\simon1.millis_counter[9] ));
 sg13g2_nor3_1 _1502_ (.A(\simon1.millis_counter[1] ),
    .B(\simon1.millis_counter[0] ),
    .C(_0839_),
    .Y(_0840_));
 sg13g2_nand2b_1 _1503_ (.Y(_0841_),
    .B(\simon1.millis_counter[3] ),
    .A_N(\simon1.millis_counter[4] ));
 sg13g2_nor3_1 _1504_ (.A(\simon1.millis_counter[7] ),
    .B(\simon1.millis_counter[6] ),
    .C(_0841_),
    .Y(_0842_));
 sg13g2_nand4_1 _1505_ (.B(\simon1.millis_counter[5] ),
    .C(_0840_),
    .A(\simon1.millis_counter[2] ),
    .Y(_0843_),
    .D(_0842_));
 sg13g2_tiehi _2615__109 (.L_HI(net109));
 sg13g2_nor2_1 _1507_ (.A(_0835_),
    .B(net43),
    .Y(_0845_));
 sg13g2_tiehi _2614__108 (.L_HI(net108));
 sg13g2_inv_1 _1509_ (.Y(_0847_),
    .A(\simon1.state[7] ));
 sg13g2_nand2b_2 _1510_ (.Y(_0848_),
    .B(_0793_),
    .A_N(net2));
 sg13g2_nor2_2 _1511_ (.A(_0847_),
    .B(_0848_),
    .Y(_0849_));
 sg13g2_a21oi_1 _1512_ (.A1(_0833_),
    .A2(_0845_),
    .Y(_0850_),
    .B1(_0849_));
 sg13g2_nor2_1 _1513_ (.A(net94),
    .B(_0850_),
    .Y(_0012_));
 sg13g2_tiehi _2613__107 (.L_HI(net107));
 sg13g2_tiehi _2609__106 (.L_HI(net106));
 sg13g2_inv_1 _1516_ (.Y(_0853_),
    .A(\simon1.state[6] ));
 sg13g2_inv_1 _1517_ (.Y(_0854_),
    .A(\simon1.millis_counter[4] ));
 sg13g2_inv_1 _1518_ (.Y(_0855_),
    .A(\simon1.millis_counter[7] ));
 sg13g2_nor4_1 _1519_ (.A(_0854_),
    .B(\simon1.millis_counter[5] ),
    .C(_0855_),
    .D(\simon1.millis_counter[6] ),
    .Y(_0856_));
 sg13g2_nand2_1 _1520_ (.Y(_0857_),
    .A(_0840_),
    .B(_0856_));
 sg13g2_nor3_1 _1521_ (.A(\simon1.millis_counter[2] ),
    .B(\simon1.millis_counter[3] ),
    .C(_0857_),
    .Y(_0858_));
 sg13g2_nor2_1 _1522_ (.A(_0853_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_tiehi _2608__105 (.L_HI(net105));
 sg13g2_tiehi _2607__104 (.L_HI(net104));
 sg13g2_o21ai_1 _1525_ (.B1(net95),
    .Y(_0862_),
    .A1(\simon1.state[2] ),
    .A2(_0859_));
 sg13g2_inv_1 _1526_ (.Y(_0011_),
    .A(_0862_));
 sg13g2_tiehi _2606__103 (.L_HI(net103));
 sg13g2_xor2_1 _1528_ (.B(net5),
    .A(net4),
    .X(_0864_));
 sg13g2_o21ai_1 _1529_ (.B1(net3),
    .Y(_0865_),
    .A1(net4),
    .A2(net5));
 sg13g2_o21ai_1 _1530_ (.B1(_0865_),
    .Y(_0866_),
    .A1(net3),
    .A2(_0864_));
 sg13g2_nand2_1 _1531_ (.Y(_0867_),
    .A(net2),
    .B(_0793_));
 sg13g2_o21ai_1 _1532_ (.B1(_0867_),
    .Y(_0868_),
    .A1(net2),
    .A2(_0866_));
 sg13g2_and2_1 _1533_ (.A(net62),
    .B(net43),
    .X(_0869_));
 sg13g2_tiehi _2605__102 (.L_HI(net102));
 sg13g2_a21oi_1 _1535_ (.A1(\simon1.state[1] ),
    .A2(_0868_),
    .Y(_0871_),
    .B1(net41));
 sg13g2_nor2_1 _1536_ (.A(net86),
    .B(_0871_),
    .Y(_0010_));
 sg13g2_tielo _2622__100 (.L_LO(net100));
 sg13g2_nor2b_1 _1538_ (.A(\simon1.millis_counter[3] ),
    .B_N(\simon1.millis_counter[2] ),
    .Y(_0873_));
 sg13g2_nand3_1 _1539_ (.B(\simon1.millis_counter[7] ),
    .C(\simon1.millis_counter[6] ),
    .A(\simon1.millis_counter[5] ),
    .Y(_0874_));
 sg13g2_inv_1 _1540_ (.Y(_0875_),
    .A(_0874_));
 sg13g2_nand4_1 _1541_ (.B(_0840_),
    .C(_0873_),
    .A(\simon1.millis_counter[4] ),
    .Y(_0876_),
    .D(_0875_));
 sg13g2_nand2_1 _1542_ (.Y(_0877_),
    .A(\simon1.state[4] ),
    .B(_0876_));
 sg13g2_o21ai_1 _1543_ (.B1(_0848_),
    .Y(_0878_),
    .A1(\simon1.state[7] ),
    .A2(\simon1.state[0] ));
 sg13g2_tielo _2620__99 (.L_LO(net99));
 sg13g2_a21oi_1 _1545_ (.A1(_0877_),
    .A2(_0878_),
    .Y(_0009_),
    .B1(net94));
 sg13g2_tielo ttsimon_98 (.L_LO(net98));
 sg13g2_buf_2 fanout97 (.A(net1),
    .X(net97));
 sg13g2_buf_2 fanout96 (.A(net1),
    .X(net96));
 sg13g2_or2_1 _1549_ (.X(_0883_),
    .B(net68),
    .A(net70));
 sg13g2_nand2b_1 _1550_ (.Y(_0884_),
    .B(\simon1.seq_counter[0] ),
    .A_N(\simon1.seq_counter[1] ));
 sg13g2_xor2_1 _1551_ (.B(\simon1.seq_counter[1] ),
    .A(_0027_),
    .X(_0885_));
 sg13g2_nand3b_1 _1552_ (.B(_0885_),
    .C(net70),
    .Y(_0886_),
    .A_N(\simon1.seq_counter[0] ));
 sg13g2_o21ai_1 _1553_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0883_),
    .A2(_0884_));
 sg13g2_o21ai_1 _1554_ (.B1(_0887_),
    .Y(_0888_),
    .A1(\simon1.seq_counter[2] ),
    .A2(_0028_));
 sg13g2_inv_1 _1555_ (.Y(_0889_),
    .A(_0028_));
 sg13g2_nand2_1 _1556_ (.Y(_0890_),
    .A(\simon1.seq_counter[2] ),
    .B(_0889_));
 sg13g2_and2_1 _1557_ (.A(\simon1.seq_counter[0] ),
    .B(\simon1.seq_counter[1] ),
    .X(_0891_));
 sg13g2_buf_2 fanout95 (.A(net96),
    .X(net95));
 sg13g2_nor2b_1 _1559_ (.A(net69),
    .B_N(_0027_),
    .Y(_0893_));
 sg13g2_nand3_1 _1560_ (.B(_0891_),
    .C(_0893_),
    .A(_0890_),
    .Y(_0894_));
 sg13g2_and2_1 _1561_ (.A(\simon1.seq_counter[2] ),
    .B(_0891_),
    .X(_0895_));
 sg13g2_buf_1 fanout94 (.A(_0796_),
    .X(net94));
 sg13g2_xor2_1 _1563_ (.B(_0895_),
    .A(_0029_),
    .X(_0897_));
 sg13g2_xor2_1 _1564_ (.B(_0030_),
    .A(\simon1.seq_counter[4] ),
    .X(_0898_));
 sg13g2_o21ai_1 _1565_ (.B1(\simon1.seq_counter[3] ),
    .Y(_0899_),
    .A1(_0029_),
    .A2(_0895_));
 sg13g2_and2_1 _1566_ (.A(_0898_),
    .B(_0899_),
    .X(_0900_));
 sg13g2_o21ai_1 _1567_ (.B1(_0900_),
    .Y(_0901_),
    .A1(\simon1.seq_counter[3] ),
    .A2(_0897_));
 sg13g2_and2_1 _1568_ (.A(\simon1.seq_counter[3] ),
    .B(_0895_),
    .X(_0902_));
 sg13g2_nand3b_1 _1569_ (.B(_0902_),
    .C(_0029_),
    .Y(_0903_),
    .A_N(_0030_));
 sg13g2_nand2_1 _1570_ (.Y(_0904_),
    .A(\simon1.seq_counter[3] ),
    .B(\simon1.seq_counter[4] ));
 sg13g2_mux2_1 _1571_ (.A0(_0889_),
    .A1(_0904_),
    .S(_0891_),
    .X(_0905_));
 sg13g2_a21oi_1 _1572_ (.A1(_0028_),
    .A2(_0891_),
    .Y(_0906_),
    .B1(\simon1.seq_counter[2] ));
 sg13g2_a21oi_1 _1573_ (.A1(\simon1.seq_counter[2] ),
    .A2(_0905_),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_a221oi_1 _1574_ (.B2(_0903_),
    .C1(_0907_),
    .B1(_0901_),
    .A1(_0888_),
    .Y(_0908_),
    .A2(_0894_));
 sg13g2_buf_1 fanout93 (.A(net94),
    .X(net93));
 sg13g2_nor3_1 _1576_ (.A(_0835_),
    .B(_0833_),
    .C(net43),
    .Y(_0910_));
 sg13g2_buf_2 fanout92 (.A(net93),
    .X(net92));
 sg13g2_inv_1 _1578_ (.Y(_0912_),
    .A(net63));
 sg13g2_buf_2 fanout91 (.A(net93),
    .X(net91));
 sg13g2_inv_1 _1580_ (.Y(_0914_),
    .A(\simon1.millis_counter[1] ));
 sg13g2_or2_1 _1581_ (.X(_0915_),
    .B(\simon1.millis_counter[8] ),
    .A(\simon1.millis_counter[9] ));
 sg13g2_nor3_1 _1582_ (.A(_0914_),
    .B(\simon1.millis_counter[0] ),
    .C(_0915_),
    .Y(_0916_));
 sg13g2_nand3_1 _1583_ (.B(_0873_),
    .C(_0916_),
    .A(_0856_),
    .Y(_0917_));
 sg13g2_buf_1 fanout90 (.A(_0796_),
    .X(net90));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_nand2_1 _1586_ (.Y(_0920_),
    .A(net59),
    .B(net57));
 sg13g2_nor3_1 _1587_ (.A(_0032_),
    .B(_0917_),
    .C(_0920_),
    .Y(_0921_));
 sg13g2_nor2_1 _1588_ (.A(_0912_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_a21oi_1 _1589_ (.A1(_0908_),
    .A2(_0910_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nor2_1 _1590_ (.A(net86),
    .B(_0923_),
    .Y(_0008_));
 sg13g2_nand2_1 _1591_ (.Y(_0924_),
    .A(\simon1.state[6] ),
    .B(_0858_));
 sg13g2_buf_2 fanout88 (.A(net90),
    .X(net88));
 sg13g2_nand2_1 _1593_ (.Y(_0926_),
    .A(net63),
    .B(_0921_));
 sg13g2_o21ai_1 _1594_ (.B1(_0926_),
    .Y(_0927_),
    .A1(_0908_),
    .A2(_0924_));
 sg13g2_inv_1 _1595_ (.Y(_0928_),
    .A(\simon1.state[4] ));
 sg13g2_nor3_1 _1596_ (.A(net94),
    .B(_0928_),
    .C(_0876_),
    .Y(_0089_));
 sg13g2_a21o_1 _1597_ (.A2(_0927_),
    .A1(net95),
    .B1(_0089_),
    .X(_0007_));
 sg13g2_inv_1 _1598_ (.Y(_0929_),
    .A(_0908_));
 sg13g2_nand2b_1 _1599_ (.Y(_0930_),
    .B(\simon1.state[1] ),
    .A_N(_0868_));
 sg13g2_o21ai_1 _1600_ (.B1(_0930_),
    .Y(_0931_),
    .A1(_0929_),
    .A2(_0924_));
 sg13g2_a21oi_1 _1601_ (.A1(_0929_),
    .A2(_0910_),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_nor2_1 _1602_ (.A(net87),
    .B(_0932_),
    .Y(_0006_));
 sg13g2_xor2_1 _1603_ (.B(net6),
    .A(\simon1.score1.active_digit ),
    .X(_0015_));
 sg13g2_inv_1 _1604_ (.Y(_0014_),
    .A(_0015_));
 sg13g2_nor4_1 _1605_ (.A(net63),
    .B(net61),
    .C(\simon1.state[6] ),
    .D(\simon1.state[4] ),
    .Y(_0933_));
 sg13g2_nand2b_1 _1606_ (.Y(_0934_),
    .B(_0933_),
    .A_N(\simon1.state[2] ));
 sg13g2_o21ai_1 _1607_ (.B1(_0033_),
    .Y(_0935_),
    .A1(\simon1.state[1] ),
    .A2(_0934_));
 sg13g2_nand2_1 _1608_ (.Y(_0936_),
    .A(_0848_),
    .B(_0935_));
 sg13g2_nand2_1 _1609_ (.Y(_0937_),
    .A(_0033_),
    .B(net95));
 sg13g2_or4_2 _1610_ (.A(\simon1.state[0] ),
    .B(_0794_),
    .C(_0937_),
    .D(_0934_),
    .X(_0938_));
 sg13g2_buf_1 fanout87 (.A(_0796_),
    .X(net87));
 sg13g2_o21ai_1 _1612_ (.B1(_0938_),
    .Y(_0940_),
    .A1(net87),
    .A2(_0936_));
 sg13g2_and2_1 _1613_ (.A(\simon1.next_random[0] ),
    .B(_0940_),
    .X(_0941_));
 sg13g2_buf_2 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_0000_));
 sg13g2_nand3_1 _1616_ (.B(_0938_),
    .C(_0936_),
    .A(net95),
    .Y(_0944_));
 sg13g2_o21ai_1 _1617_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0893_),
    .A2(_0938_));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_0000_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_0001_));
 sg13g2_nor3_1 _1620_ (.A(net67),
    .B(net66),
    .C(\simon1.seq_length[4] ),
    .Y(_0948_));
 sg13g2_nor4_2 _1621_ (.A(\simon1.state[0] ),
    .B(_0794_),
    .C(_0937_),
    .Y(_0949_),
    .D(_0934_));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_0001_));
 sg13g2_nand2b_1 _1623_ (.Y(_0951_),
    .B(_0949_),
    .A_N(_0948_));
 sg13g2_nor2b_1 _1624_ (.A(_0945_),
    .B_N(_0951_),
    .Y(_0952_));
 sg13g2_mux2_1 _1625_ (.A0(\simon1.seq[0][0] ),
    .A1(net32),
    .S(_0952_),
    .X(_0038_));
 sg13g2_and2_1 _1626_ (.A(\simon1.next_random[1] ),
    .B(_0940_),
    .X(_0953_));
 sg13g2_buf_2 fanout81 (.A(\simon1.play1.freq[5] ),
    .X(net81));
 sg13g2_buf_1 fanout80 (.A(\simon1.play1.freq[6] ),
    .X(net80));
 sg13g2_nor2_1 _1629_ (.A(net67),
    .B(\simon1.seq_length[4] ),
    .Y(_0956_));
 sg13g2_nand3_1 _1630_ (.B(_0949_),
    .C(_0956_),
    .A(net66),
    .Y(_0957_));
 sg13g2_nor2_1 _1631_ (.A(_0945_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_mux2_1 _1632_ (.A0(\simon1.seq[8][1] ),
    .A1(net28),
    .S(_0958_),
    .X(_0039_));
 sg13g2_nand2_1 _1633_ (.Y(_0959_),
    .A(net67),
    .B(net42));
 sg13g2_or2_1 _1634_ (.X(_0960_),
    .B(_0959_),
    .A(\simon1.seq_length[4] ));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_1 fanout78 (.A(\simon1.play1.freq[8] ),
    .X(net78));
 sg13g2_nor2_1 _1637_ (.A(net69),
    .B(net68),
    .Y(_0963_));
 sg13g2_nand2_1 _1638_ (.Y(_0964_),
    .A(net65),
    .B(_0963_));
 sg13g2_nor2_1 _1639_ (.A(_0960_),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_mux2_1 _1640_ (.A0(\simon1.seq[14][1] ),
    .A1(net28),
    .S(_0965_),
    .X(_0040_));
 sg13g2_and3_1 _1641_ (.X(_0966_),
    .A(net69),
    .B(net68),
    .C(net42));
 sg13g2_nand2_1 _1642_ (.Y(_0967_),
    .A(net66),
    .B(_0966_));
 sg13g2_nor2_1 _1643_ (.A(_0960_),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_mux2_1 _1644_ (.A0(\simon1.seq[13][1] ),
    .A1(net28),
    .S(_0968_),
    .X(_0041_));
 sg13g2_inv_1 _1645_ (.Y(_0969_),
    .A(_0945_));
 sg13g2_nand2_1 _1646_ (.Y(_0970_),
    .A(net65),
    .B(_0969_));
 sg13g2_nor2_1 _1647_ (.A(_0960_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_mux2_1 _1648_ (.A0(\simon1.seq[12][1] ),
    .A1(net28),
    .S(_0971_),
    .X(_0042_));
 sg13g2_buf_2 fanout77 (.A(net78),
    .X(net77));
 sg13g2_nor2b_1 _1650_ (.A(net68),
    .B_N(net69),
    .Y(_0973_));
 sg13g2_nand3_1 _1651_ (.B(_0948_),
    .C(_0973_),
    .A(net42),
    .Y(_0974_));
 sg13g2_mux2_1 _1652_ (.A0(net32),
    .A1(\simon1.seq[3][0] ),
    .S(_0974_),
    .X(_0043_));
 sg13g2_nand3_1 _1653_ (.B(\simon1.seq_length[4] ),
    .C(net42),
    .A(net67),
    .Y(_0975_));
 sg13g2_nand2_1 _1654_ (.Y(_0976_),
    .A(net65),
    .B(_0973_));
 sg13g2_or2_1 _1655_ (.X(_0977_),
    .B(_0976_),
    .A(_0975_));
 sg13g2_mux2_1 _1656_ (.A0(net34),
    .A1(\simon1.seq[31][0] ),
    .S(_0977_),
    .X(_0044_));
 sg13g2_nand3_1 _1657_ (.B(net42),
    .C(_0948_),
    .A(_0963_),
    .Y(_0978_));
 sg13g2_mux2_1 _1658_ (.A0(net32),
    .A1(\simon1.seq[2][0] ),
    .S(_0978_),
    .X(_0045_));
 sg13g2_nor2_1 _1659_ (.A(_0967_),
    .B(_0975_),
    .Y(_0979_));
 sg13g2_mux2_1 _1660_ (.A0(\simon1.seq[29][0] ),
    .A1(net30),
    .S(_0979_),
    .X(_0046_));
 sg13g2_nor2_1 _1661_ (.A(_0970_),
    .B(_0975_),
    .Y(_0980_));
 sg13g2_mux2_1 _1662_ (.A0(\simon1.seq[28][0] ),
    .A1(net30),
    .S(_0980_),
    .X(_0047_));
 sg13g2_nand3b_1 _1663_ (.B(\simon1.seq_length[4] ),
    .C(net42),
    .Y(_0981_),
    .A_N(net67));
 sg13g2_buf_2 fanout76 (.A(\simon1.play1.tick_counter[11] ),
    .X(net76));
 sg13g2_nor2_1 _1665_ (.A(_0976_),
    .B(_0981_),
    .Y(_0983_));
 sg13g2_mux2_1 _1666_ (.A0(\simon1.seq[27][0] ),
    .A1(net30),
    .S(_0983_),
    .X(_0048_));
 sg13g2_nor2_1 _1667_ (.A(_0964_),
    .B(_0981_),
    .Y(_0984_));
 sg13g2_mux2_1 _1668_ (.A0(\simon1.seq[26][0] ),
    .A1(net30),
    .S(_0984_),
    .X(_0049_));
 sg13g2_or2_1 _1669_ (.X(_0985_),
    .B(_0981_),
    .A(_0967_));
 sg13g2_mux2_1 _1670_ (.A0(net30),
    .A1(\simon1.seq[25][0] ),
    .S(_0985_),
    .X(_0050_));
 sg13g2_or2_1 _1671_ (.X(_0986_),
    .B(_0981_),
    .A(_0970_));
 sg13g2_mux2_1 _1672_ (.A0(net30),
    .A1(\simon1.seq[24][0] ),
    .S(_0986_),
    .X(_0051_));
 sg13g2_and3_1 _1673_ (.X(_0987_),
    .A(net67),
    .B(\simon1.seq_length[4] ),
    .C(net42));
 sg13g2_buf_2 fanout75 (.A(\simon1.play1.tick_counter[12] ),
    .X(net75));
 sg13g2_buf_2 fanout74 (.A(\simon1.play1.tick_counter[27] ),
    .X(net74));
 sg13g2_nand2b_1 _1676_ (.Y(_0990_),
    .B(net69),
    .A_N(net68));
 sg13g2_nor2_1 _1677_ (.A(net65),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_nand2_1 _1678_ (.Y(_0992_),
    .A(_0987_),
    .B(_0991_));
 sg13g2_mux2_1 _1679_ (.A0(net31),
    .A1(\simon1.seq[23][0] ),
    .S(_0992_),
    .X(_0052_));
 sg13g2_nor3_2 _1680_ (.A(net69),
    .B(net68),
    .C(net65),
    .Y(_0993_));
 sg13g2_nand2_1 _1681_ (.Y(_0994_),
    .A(_0987_),
    .B(_0993_));
 sg13g2_mux2_1 _1682_ (.A0(net31),
    .A1(\simon1.seq[22][0] ),
    .S(_0994_),
    .X(_0053_));
 sg13g2_nor3_1 _1683_ (.A(_0938_),
    .B(_0957_),
    .C(_0990_),
    .Y(_0995_));
 sg13g2_mux2_1 _1684_ (.A0(\simon1.seq[11][1] ),
    .A1(net27),
    .S(_0995_),
    .X(_0054_));
 sg13g2_nand3_1 _1685_ (.B(net68),
    .C(net42),
    .A(net69),
    .Y(_0996_));
 sg13g2_nor2_1 _1686_ (.A(net65),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_nand2_1 _1687_ (.Y(_0998_),
    .A(_0987_),
    .B(_0997_));
 sg13g2_mux2_1 _1688_ (.A0(net31),
    .A1(\simon1.seq[21][0] ),
    .S(_0998_),
    .X(_0055_));
 sg13g2_nand2_1 _1689_ (.Y(_0999_),
    .A(_0951_),
    .B(_0966_));
 sg13g2_mux2_1 _1690_ (.A0(net32),
    .A1(\simon1.seq[1][0] ),
    .S(_0999_),
    .X(_0056_));
 sg13g2_nand2b_1 _1691_ (.Y(_1000_),
    .B(_0991_),
    .A_N(_0981_));
 sg13g2_mux2_1 _1692_ (.A0(net31),
    .A1(\simon1.seq[19][0] ),
    .S(_1000_),
    .X(_0057_));
 sg13g2_nand2b_1 _1693_ (.Y(_1001_),
    .B(_0993_),
    .A_N(_0981_));
 sg13g2_mux2_1 _1694_ (.A0(net31),
    .A1(\simon1.seq[18][0] ),
    .S(_1001_),
    .X(_0058_));
 sg13g2_buf_2 fanout73 (.A(\simon1.play1.tick_counter[5] ),
    .X(net73));
 sg13g2_nor3_1 _1696_ (.A(net65),
    .B(_0996_),
    .C(_0981_),
    .Y(_1003_));
 sg13g2_mux2_1 _1697_ (.A0(\simon1.seq[17][0] ),
    .A1(net30),
    .S(_1003_),
    .X(_0059_));
 sg13g2_or2_1 _1698_ (.X(_1004_),
    .B(_0945_),
    .A(net65));
 sg13g2_nor2_1 _1699_ (.A(_0981_),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_mux2_1 _1700_ (.A0(\simon1.seq[16][0] ),
    .A1(net31),
    .S(_1005_),
    .X(_0060_));
 sg13g2_nor2_1 _1701_ (.A(_0960_),
    .B(_0976_),
    .Y(_1006_));
 sg13g2_mux2_1 _1702_ (.A0(\simon1.seq[15][0] ),
    .A1(net33),
    .S(_1006_),
    .X(_0061_));
 sg13g2_mux2_1 _1703_ (.A0(\simon1.seq[14][0] ),
    .A1(net33),
    .S(_0965_),
    .X(_0062_));
 sg13g2_mux2_1 _1704_ (.A0(\simon1.seq[13][0] ),
    .A1(net33),
    .S(_0968_),
    .X(_0063_));
 sg13g2_buf_2 fanout72 (.A(\simon1.play1.tick_counter[8] ),
    .X(net72));
 sg13g2_nor4_2 _1706_ (.A(net69),
    .B(net68),
    .C(_0938_),
    .Y(_1008_),
    .D(_0957_));
 sg13g2_mux2_1 _1707_ (.A0(\simon1.seq[10][1] ),
    .A1(net28),
    .S(_1008_),
    .X(_0064_));
 sg13g2_mux2_1 _1708_ (.A0(\simon1.seq[12][0] ),
    .A1(net33),
    .S(_0971_),
    .X(_0065_));
 sg13g2_mux2_1 _1709_ (.A0(\simon1.seq[11][0] ),
    .A1(net32),
    .S(_0995_),
    .X(_0066_));
 sg13g2_nor2_1 _1710_ (.A(_0957_),
    .B(_0996_),
    .Y(_1009_));
 sg13g2_mux2_1 _1711_ (.A0(\simon1.seq[9][1] ),
    .A1(net28),
    .S(_1009_),
    .X(_0067_));
 sg13g2_mux2_1 _1712_ (.A0(\simon1.seq[9][0] ),
    .A1(net33),
    .S(_1009_),
    .X(_0068_));
 sg13g2_buf_2 fanout71 (.A(\simon1.score1.active_digit ),
    .X(net71));
 sg13g2_nor2_1 _1714_ (.A(\simon1.seq_length[4] ),
    .B(_0959_),
    .Y(_1011_));
 sg13g2_nand2_1 _1715_ (.Y(_1012_),
    .A(_1011_),
    .B(_0991_));
 sg13g2_mux2_1 _1716_ (.A0(net27),
    .A1(\simon1.seq[7][1] ),
    .S(_1012_),
    .X(_0069_));
 sg13g2_nand2_1 _1717_ (.Y(_1013_),
    .A(_1011_),
    .B(_0993_));
 sg13g2_mux2_1 _1718_ (.A0(net27),
    .A1(\simon1.seq[6][1] ),
    .S(_1013_),
    .X(_0070_));
 sg13g2_nand2_1 _1719_ (.Y(_1014_),
    .A(_1011_),
    .B(_0997_));
 sg13g2_mux2_1 _1720_ (.A0(net27),
    .A1(\simon1.seq[5][1] ),
    .S(_1014_),
    .X(_0071_));
 sg13g2_mux2_1 _1721_ (.A0(\simon1.seq[8][0] ),
    .A1(net33),
    .S(_0958_),
    .X(_0072_));
 sg13g2_mux2_1 _1722_ (.A0(net32),
    .A1(\simon1.seq[7][0] ),
    .S(_1012_),
    .X(_0073_));
 sg13g2_mux2_1 _1723_ (.A0(net32),
    .A1(\simon1.seq[6][0] ),
    .S(_1013_),
    .X(_0074_));
 sg13g2_mux2_1 _1724_ (.A0(net32),
    .A1(\simon1.seq[5][0] ),
    .S(_1014_),
    .X(_0075_));
 sg13g2_nor2_1 _1725_ (.A(_0960_),
    .B(_1004_),
    .Y(_1015_));
 sg13g2_mux2_1 _1726_ (.A0(\simon1.seq[4][1] ),
    .A1(net26),
    .S(_1015_),
    .X(_0076_));
 sg13g2_mux2_1 _1727_ (.A0(net29),
    .A1(\simon1.seq[31][1] ),
    .S(_0977_),
    .X(_0077_));
 sg13g2_mux2_1 _1728_ (.A0(net27),
    .A1(\simon1.seq[3][1] ),
    .S(_0974_),
    .X(_0078_));
 sg13g2_mux2_1 _1729_ (.A0(\simon1.seq[4][0] ),
    .A1(net31),
    .S(_1015_),
    .X(_0079_));
 sg13g2_nand2b_1 _1730_ (.Y(_1016_),
    .B(_0987_),
    .A_N(_0964_));
 sg13g2_mux2_1 _1731_ (.A0(net30),
    .A1(\simon1.seq[30][0] ),
    .S(_1016_),
    .X(_0080_));
 sg13g2_mux2_1 _1732_ (.A0(net25),
    .A1(\simon1.seq[30][1] ),
    .S(_1016_),
    .X(_0087_));
 sg13g2_mux2_1 _1733_ (.A0(net27),
    .A1(\simon1.seq[2][1] ),
    .S(_0978_),
    .X(_0088_));
 sg13g2_mux2_1 _1734_ (.A0(\simon1.seq[28][1] ),
    .A1(net25),
    .S(_0980_),
    .X(_0131_));
 sg13g2_nor2_1 _1735_ (.A(net3),
    .B(net5),
    .Y(_1017_));
 sg13g2_nand2_1 _1736_ (.Y(_1018_),
    .A(net97),
    .B(\simon1.state[1] ));
 sg13g2_nand2b_1 _1737_ (.Y(_1019_),
    .B(net4),
    .A_N(net2));
 sg13g2_o21ai_1 _1738_ (.B1(\simon1.user_input[0] ),
    .Y(_1020_),
    .A1(_1018_),
    .A2(_1019_));
 sg13g2_nor2_1 _1739_ (.A(net4),
    .B(_1018_),
    .Y(_1021_));
 sg13g2_inv_1 _1740_ (.Y(_1022_),
    .A(\simon1.user_input[0] ));
 sg13g2_a21o_1 _1741_ (.A2(_1021_),
    .A1(_1017_),
    .B1(_1022_),
    .X(_1023_));
 sg13g2_nand2_1 _1742_ (.Y(_1024_),
    .A(net3),
    .B(net5));
 sg13g2_a21oi_1 _1743_ (.A1(_1021_),
    .A2(_1024_),
    .Y(_1025_),
    .B1(\simon1.user_input[0] ));
 sg13g2_a221oi_1 _1744_ (.B2(net2),
    .C1(_1025_),
    .B1(_1023_),
    .A1(_1017_),
    .Y(_0134_),
    .A2(_1020_));
 sg13g2_inv_1 _1745_ (.Y(_1026_),
    .A(\simon1.user_input[1] ));
 sg13g2_nand2b_1 _1746_ (.Y(_1027_),
    .B(_0864_),
    .A_N(_1018_));
 sg13g2_nand2b_1 _1747_ (.Y(_1028_),
    .B(_1021_),
    .A_N(net5));
 sg13g2_nand3_1 _1748_ (.B(net2),
    .C(net3),
    .A(\simon1.user_input[1] ),
    .Y(_1029_));
 sg13g2_o21ai_1 _1749_ (.B1(_1029_),
    .Y(_1030_),
    .A1(net2),
    .A2(net3));
 sg13g2_a21oi_1 _1750_ (.A1(\simon1.user_input[1] ),
    .A2(_1028_),
    .Y(_1031_),
    .B1(_1030_));
 sg13g2_a21oi_1 _1751_ (.A1(_1026_),
    .A2(_1027_),
    .Y(_0135_),
    .B1(_1031_));
 sg13g2_buf_2 fanout70 (.A(\simon1.seq_length[0] ),
    .X(net70));
 sg13g2_inv_1 _1753_ (.Y(_1033_),
    .A(_0034_));
 sg13g2_inv_1 _1754_ (.Y(_1034_),
    .A(net58));
 sg13g2_nand2_1 _1755_ (.Y(_1035_),
    .A(net55),
    .B(_1034_));
 sg13g2_a21oi_1 _1756_ (.A1(net60),
    .A2(_1033_),
    .Y(_1036_),
    .B1(_1035_));
 sg13g2_nor3_1 _1757_ (.A(_0847_),
    .B(_0032_),
    .C(_1036_),
    .Y(_1037_));
 sg13g2_nor2_2 _1758_ (.A(net60),
    .B(net58),
    .Y(_1038_));
 sg13g2_and2_1 _1759_ (.A(net56),
    .B(_1038_),
    .X(_1039_));
 sg13g2_buf_2 fanout69 (.A(\simon1.seq_length[0] ),
    .X(net69));
 sg13g2_o21ai_1 _1761_ (.B1(_0843_),
    .Y(_1041_),
    .A1(_0033_),
    .A2(_1039_));
 sg13g2_o21ai_1 _1762_ (.B1(_1041_),
    .Y(_1042_),
    .A1(net43),
    .A2(_1037_));
 sg13g2_nor2_1 _1763_ (.A(net63),
    .B(\simon1.state[4] ),
    .Y(_1043_));
 sg13g2_a21oi_1 _1764_ (.A1(_0033_),
    .A2(_1043_),
    .Y(_1044_),
    .B1(net86));
 sg13g2_and2_1 _1765_ (.A(net63),
    .B(_0917_),
    .X(_1045_));
 sg13g2_buf_2 fanout68 (.A(_0027_),
    .X(net68));
 sg13g2_nand2_2 _1767_ (.Y(_1047_),
    .A(net56),
    .B(_1038_));
 sg13g2_nand2_1 _1768_ (.Y(_1048_),
    .A(\simon1.millis_counter[9] ),
    .B(\simon1.millis_counter[8] ));
 sg13g2_nor3_1 _1769_ (.A(_0841_),
    .B(_0874_),
    .C(_1048_),
    .Y(_1049_));
 sg13g2_nor3_1 _1770_ (.A(\simon1.millis_counter[1] ),
    .B(\simon1.millis_counter[0] ),
    .C(\simon1.millis_counter[2] ),
    .Y(_1050_));
 sg13g2_and2_1 _1771_ (.A(_1049_),
    .B(_1050_),
    .X(_1051_));
 sg13g2_buf_2 fanout67 (.A(\simon1.seq_length[2] ),
    .X(net67));
 sg13g2_nor3_1 _1773_ (.A(_0847_),
    .B(_1047_),
    .C(_1051_),
    .Y(_1053_));
 sg13g2_nor2_1 _1774_ (.A(_1045_),
    .B(_1053_),
    .Y(_1054_));
 sg13g2_nand3_1 _1775_ (.B(_1044_),
    .C(_1054_),
    .A(_1042_),
    .Y(_1055_));
 sg13g2_buf_1 fanout66 (.A(\simon1.seq_length[3] ),
    .X(net66));
 sg13g2_nor2_1 _1777_ (.A(\simon1.state[7] ),
    .B(net63),
    .Y(_1057_));
 sg13g2_nor3_1 _1778_ (.A(net59),
    .B(_1055_),
    .C(_1057_),
    .Y(_1058_));
 sg13g2_a21o_1 _1779_ (.A2(_1055_),
    .A1(net59),
    .B1(_1058_),
    .X(_0138_));
 sg13g2_inv_1 _1780_ (.Y(_1059_),
    .A(net59));
 sg13g2_inv_1 _1781_ (.Y(_1060_),
    .A(_0033_));
 sg13g2_nand2_1 _1782_ (.Y(_1061_),
    .A(net55),
    .B(_1060_));
 sg13g2_a21oi_1 _1783_ (.A1(_1059_),
    .A2(_1061_),
    .Y(_1062_),
    .B1(_1055_));
 sg13g2_nor2_1 _1784_ (.A(net57),
    .B(_1062_),
    .Y(_1063_));
 sg13g2_a21oi_1 _1785_ (.A1(\simon1.state[7] ),
    .A2(_1060_),
    .Y(_1064_),
    .B1(net63));
 sg13g2_a21oi_1 _1786_ (.A1(net59),
    .A2(net57),
    .Y(_1065_),
    .B1(_1064_));
 sg13g2_nor2_1 _1787_ (.A(_1055_),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nor2_1 _1788_ (.A(_1063_),
    .B(_1066_),
    .Y(_0139_));
 sg13g2_o21ai_1 _1789_ (.B1(_0032_),
    .Y(_1067_),
    .A1(net57),
    .A2(_1061_));
 sg13g2_nand2_1 _1790_ (.Y(_1068_),
    .A(_0032_),
    .B(_0920_));
 sg13g2_inv_1 _1791_ (.Y(_1069_),
    .A(_0032_));
 sg13g2_nand2_1 _1792_ (.Y(_1070_),
    .A(net57),
    .B(_1069_));
 sg13g2_a22oi_1 _1793_ (.Y(_1071_),
    .B1(_1068_),
    .B2(_1070_),
    .A2(_1067_),
    .A1(_1059_));
 sg13g2_nor3_1 _1794_ (.A(_1055_),
    .B(_1064_),
    .C(_1071_),
    .Y(_1072_));
 sg13g2_a21o_1 _1795_ (.A2(_1055_),
    .A1(net55),
    .B1(_1072_),
    .X(_0140_));
 sg13g2_mux2_1 _1796_ (.A0(\simon1.seq[27][1] ),
    .A1(net25),
    .S(_0983_),
    .X(_0186_));
 sg13g2_mux2_1 _1797_ (.A0(net26),
    .A1(\simon1.seq[18][1] ),
    .S(_1001_),
    .X(_0187_));
 sg13g2_mux2_1 _1798_ (.A0(\simon1.seq[26][1] ),
    .A1(net25),
    .S(_0984_),
    .X(_0188_));
 sg13g2_mux2_1 _1799_ (.A0(net25),
    .A1(\simon1.seq[25][1] ),
    .S(_0985_),
    .X(_0189_));
 sg13g2_mux2_1 _1800_ (.A0(net26),
    .A1(\simon1.seq[22][1] ),
    .S(_0994_),
    .X(_0190_));
 sg13g2_mux2_1 _1801_ (.A0(net26),
    .A1(\simon1.seq[23][1] ),
    .S(_0992_),
    .X(_0191_));
 sg13g2_nor2_1 _1802_ (.A(_0975_),
    .B(_1004_),
    .Y(_1073_));
 sg13g2_mux2_1 _1803_ (.A0(\simon1.seq[20][1] ),
    .A1(net26),
    .S(_1073_),
    .X(_0192_));
 sg13g2_mux2_1 _1804_ (.A0(net26),
    .A1(\simon1.seq[21][1] ),
    .S(_0998_),
    .X(_0193_));
 sg13g2_mux2_1 _1805_ (.A0(net25),
    .A1(\simon1.seq[24][1] ),
    .S(_0986_),
    .X(_0194_));
 sg13g2_mux2_1 _1806_ (.A0(net26),
    .A1(\simon1.seq[19][1] ),
    .S(_1000_),
    .X(_0195_));
 sg13g2_mux2_1 _1807_ (.A0(\simon1.seq[17][1] ),
    .A1(net25),
    .S(_1003_),
    .X(_0196_));
 sg13g2_mux2_1 _1808_ (.A0(\simon1.seq[10][0] ),
    .A1(net33),
    .S(_1008_),
    .X(_0197_));
 sg13g2_mux2_1 _1809_ (.A0(\simon1.seq[16][1] ),
    .A1(net26),
    .S(_1005_),
    .X(_0198_));
 sg13g2_mux2_1 _1810_ (.A0(\simon1.seq[20][0] ),
    .A1(net31),
    .S(_1073_),
    .X(_0199_));
 sg13g2_mux2_1 _1811_ (.A0(net27),
    .A1(\simon1.seq[1][1] ),
    .S(_0999_),
    .X(_0200_));
 sg13g2_mux2_1 _1812_ (.A0(\simon1.seq[15][1] ),
    .A1(net28),
    .S(_1006_),
    .X(_0201_));
 sg13g2_mux2_1 _1813_ (.A0(\simon1.seq[29][1] ),
    .A1(net25),
    .S(_0979_),
    .X(_0202_));
 sg13g2_mux2_1 _1814_ (.A0(\simon1.seq[0][1] ),
    .A1(net27),
    .S(_0952_),
    .X(_0203_));
 sg13g2_inv_1 _1815_ (.Y(_1074_),
    .A(_0016_));
 sg13g2_nand2b_1 _1816_ (.Y(_1075_),
    .B(net97),
    .A_N(\simon1.score_rst ));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_nor2_1 _1818_ (.A(_1074_),
    .B(_1075_),
    .Y(_0081_));
 sg13g2_xnor2_1 _1819_ (.Y(_1077_),
    .A(\simon1.score1.ones[0] ),
    .B(\simon1.score1.inc ));
 sg13g2_nor2_1 _1820_ (.A(net54),
    .B(_1077_),
    .Y(_0090_));
 sg13g2_nand2_2 _1821_ (.Y(_1078_),
    .A(\simon1.score1.ones[0] ),
    .B(\simon1.score1.inc ));
 sg13g2_nor2_1 _1822_ (.A(\simon1.score1.ones[2] ),
    .B(_0760_),
    .Y(_1079_));
 sg13g2_nor3_1 _1823_ (.A(\simon1.score1.ones[1] ),
    .B(_1078_),
    .C(_1079_),
    .Y(_1080_));
 sg13g2_a21oi_1 _1824_ (.A1(\simon1.score1.ones[1] ),
    .A2(_1078_),
    .Y(_1081_),
    .B1(_1080_));
 sg13g2_nor2_1 _1825_ (.A(net54),
    .B(_1081_),
    .Y(_0091_));
 sg13g2_inv_1 _1826_ (.Y(_1082_),
    .A(\simon1.score1.ones[2] ));
 sg13g2_nand3_1 _1827_ (.B(\simon1.score1.ones[1] ),
    .C(\simon1.score1.inc ),
    .A(\simon1.score1.ones[0] ),
    .Y(_1083_));
 sg13g2_xnor2_1 _1828_ (.Y(_1084_),
    .A(_1082_),
    .B(_1083_));
 sg13g2_nor2_1 _1829_ (.A(net54),
    .B(_1084_),
    .Y(_0092_));
 sg13g2_nor2_1 _1830_ (.A(\simon1.score1.ones[1] ),
    .B(_1082_),
    .Y(_1085_));
 sg13g2_o21ai_1 _1831_ (.B1(\simon1.score1.ones[3] ),
    .Y(_1086_),
    .A1(_1078_),
    .A2(_1085_));
 sg13g2_nor3_1 _1832_ (.A(_1082_),
    .B(\simon1.score1.ones[3] ),
    .C(_1078_),
    .Y(_1087_));
 sg13g2_o21ai_1 _1833_ (.B1(\simon1.score1.ones[1] ),
    .Y(_1088_),
    .A1(_1079_),
    .A2(_1087_));
 sg13g2_a21oi_1 _1834_ (.A1(_1086_),
    .A2(_1088_),
    .Y(_0093_),
    .B1(net54));
 sg13g2_nor4_2 _1835_ (.A(\simon1.score1.ones[1] ),
    .B(\simon1.score1.ones[2] ),
    .C(_0760_),
    .Y(_1089_),
    .D(_1078_));
 sg13g2_xnor2_1 _1836_ (.Y(_1090_),
    .A(\simon1.score1.tens[0] ),
    .B(_1089_));
 sg13g2_nor2_1 _1837_ (.A(net54),
    .B(_1090_),
    .Y(_0094_));
 sg13g2_nand2_1 _1838_ (.Y(_1091_),
    .A(\simon1.score1.tens[0] ),
    .B(_1089_));
 sg13g2_nor2b_1 _1839_ (.A(\simon1.score1.tens[2] ),
    .B_N(\simon1.score1.tens[3] ),
    .Y(_1092_));
 sg13g2_nor3_1 _1840_ (.A(\simon1.score1.tens[1] ),
    .B(_1091_),
    .C(_1092_),
    .Y(_1093_));
 sg13g2_a21oi_1 _1841_ (.A1(\simon1.score1.tens[1] ),
    .A2(_1091_),
    .Y(_1094_),
    .B1(_1093_));
 sg13g2_nor2_1 _1842_ (.A(net54),
    .B(_1094_),
    .Y(_0095_));
 sg13g2_nand3_1 _1843_ (.B(\simon1.score1.tens[1] ),
    .C(_1089_),
    .A(\simon1.score1.tens[0] ),
    .Y(_1095_));
 sg13g2_xnor2_1 _1844_ (.Y(_1096_),
    .A(_0755_),
    .B(_1095_));
 sg13g2_nor2_1 _1845_ (.A(net54),
    .B(_1096_),
    .Y(_0096_));
 sg13g2_nor2_1 _1846_ (.A(\simon1.score1.tens[1] ),
    .B(_0755_),
    .Y(_1097_));
 sg13g2_o21ai_1 _1847_ (.B1(\simon1.score1.tens[3] ),
    .Y(_1098_),
    .A1(_1091_),
    .A2(_1097_));
 sg13g2_nor3_1 _1848_ (.A(_0755_),
    .B(\simon1.score1.tens[3] ),
    .C(_1091_),
    .Y(_1099_));
 sg13g2_o21ai_1 _1849_ (.B1(\simon1.score1.tens[1] ),
    .Y(_1100_),
    .A1(_1092_),
    .A2(_1099_));
 sg13g2_a21oi_1 _1850_ (.A1(_1098_),
    .A2(_1100_),
    .Y(_0097_),
    .B1(net54));
 sg13g2_buf_1 fanout64 (.A(\simon1.state[3] ),
    .X(net64));
 sg13g2_and2_1 _1852_ (.A(\simon1.play1.tick_counter[14] ),
    .B(\simon1.play1.tick_counter[13] ),
    .X(_1102_));
 sg13g2_buf_2 fanout63 (.A(\simon1.state[3] ),
    .X(net63));
 sg13g2_buf_2 fanout62 (.A(\simon1.state[5] ),
    .X(net62));
 sg13g2_buf_2 fanout61 (.A(net62),
    .X(net61));
 sg13g2_nand2_1 _1856_ (.Y(_1106_),
    .A(\simon1.play1.tick_counter[7] ),
    .B(net72));
 sg13g2_buf_1 fanout60 (.A(\simon1.tone_sequence_counter[0] ),
    .X(net60));
 sg13g2_buf_2 fanout59 (.A(\simon1.tone_sequence_counter[0] ),
    .X(net59));
 sg13g2_buf_1 fanout58 (.A(\simon1.tone_sequence_counter[1] ),
    .X(net58));
 sg13g2_buf_2 fanout57 (.A(net58),
    .X(net57));
 sg13g2_o21ai_1 _1861_ (.B1(net73),
    .Y(_1111_),
    .A1(\simon1.play1.tick_counter[3] ),
    .A2(\simon1.play1.tick_counter[4] ));
 sg13g2_nor2b_1 _1862_ (.A(\simon1.play1.tick_counter[6] ),
    .B_N(_1111_),
    .Y(_1112_));
 sg13g2_buf_1 fanout56 (.A(\simon1.tone_sequence_counter[2] ),
    .X(net56));
 sg13g2_buf_2 fanout55 (.A(\simon1.tone_sequence_counter[2] ),
    .X(net55));
 sg13g2_buf_2 fanout54 (.A(_1075_),
    .X(net54));
 sg13g2_buf_2 fanout53 (.A(_0608_),
    .X(net53));
 sg13g2_nor4_1 _1867_ (.A(net75),
    .B(net76),
    .C(\simon1.play1.tick_counter[10] ),
    .D(\simon1.play1.tick_counter[9] ),
    .Y(_1117_));
 sg13g2_o21ai_1 _1868_ (.B1(_1117_),
    .Y(_1118_),
    .A1(_1106_),
    .A2(_1112_));
 sg13g2_nand2_1 _1869_ (.Y(_1119_),
    .A(_1102_),
    .B(_1118_));
 sg13g2_buf_2 fanout52 (.A(_1150_),
    .X(net52));
 sg13g2_nor3_1 _1871_ (.A(\simon1.play1.tick_counter[15] ),
    .B(\simon1.play1.tick_counter[31] ),
    .C(\simon1.play1.tick_counter[16] ),
    .Y(_1121_));
 sg13g2_buf_1 fanout51 (.A(_1232_),
    .X(net51));
 sg13g2_buf_2 fanout50 (.A(_1232_),
    .X(net50));
 sg13g2_nor4_1 _1874_ (.A(\simon1.play1.tick_counter[26] ),
    .B(\simon1.play1.tick_counter[25] ),
    .C(\simon1.play1.tick_counter[24] ),
    .D(\simon1.play1.tick_counter[23] ),
    .Y(_1124_));
 sg13g2_buf_1 fanout49 (.A(_1232_),
    .X(net49));
 sg13g2_buf_2 fanout48 (.A(net49),
    .X(net48));
 sg13g2_nor4_1 _1877_ (.A(\simon1.play1.tick_counter[30] ),
    .B(\simon1.play1.tick_counter[21] ),
    .C(\simon1.play1.tick_counter[20] ),
    .D(\simon1.play1.tick_counter[17] ),
    .Y(_1127_));
 sg13g2_nand3_1 _1878_ (.B(_1124_),
    .C(_1127_),
    .A(_1121_),
    .Y(_1128_));
 sg13g2_or2_1 _1879_ (.X(_1129_),
    .B(\simon1.play1.tick_counter[28] ),
    .A(\simon1.play1.tick_counter[29] ));
 sg13g2_buf_1 fanout47 (.A(net49),
    .X(net47));
 sg13g2_buf_2 fanout46 (.A(net49),
    .X(net46));
 sg13g2_or4_1 _1882_ (.A(net74),
    .B(\simon1.play1.tick_counter[22] ),
    .C(\simon1.play1.tick_counter[19] ),
    .D(\simon1.play1.tick_counter[18] ),
    .X(_1132_));
 sg13g2_nor3_1 _1883_ (.A(_1128_),
    .B(_1129_),
    .C(_1132_),
    .Y(_1133_));
 sg13g2_and2_2 _1884_ (.A(_1119_),
    .B(_1133_),
    .X(_1134_));
 sg13g2_buf_2 fanout45 (.A(_0440_),
    .X(net45));
 sg13g2_mux2_1 _1886_ (.A0(_0013_),
    .A1(net18),
    .S(_1134_),
    .X(_1136_));
 sg13g2_buf_2 fanout44 (.A(_0816_),
    .X(net44));
 sg13g2_buf_2 fanout43 (.A(_0843_),
    .X(net43));
 sg13g2_nor2_1 _1889_ (.A(net81),
    .B(\simon1.play1.freq[4] ),
    .Y(_1139_));
 sg13g2_buf_2 fanout42 (.A(_0949_),
    .X(net42));
 sg13g2_buf_2 fanout41 (.A(_0869_),
    .X(net41));
 sg13g2_nor2_1 _1892_ (.A(\simon1.play1.freq[9] ),
    .B(net78),
    .Y(_1142_));
 sg13g2_buf_2 fanout40 (.A(_1161_),
    .X(net40));
 sg13g2_buf_2 fanout39 (.A(net40),
    .X(net39));
 sg13g2_nor2_1 _1895_ (.A(\simon1.play1.freq[7] ),
    .B(net80),
    .Y(_1145_));
 sg13g2_buf_2 fanout38 (.A(_0358_),
    .X(net38));
 sg13g2_buf_1 fanout37 (.A(_0358_),
    .X(net37));
 sg13g2_buf_1 fanout36 (.A(net37),
    .X(net36));
 sg13g2_nor4_1 _1899_ (.A(\simon1.play1.freq[0] ),
    .B(\simon1.play1.freq[1] ),
    .C(\simon1.play1.freq[3] ),
    .D(\simon1.play1.freq[2] ),
    .Y(_1149_));
 sg13g2_nand4_1 _1900_ (.B(_1142_),
    .C(_1145_),
    .A(_1139_),
    .Y(_1150_),
    .D(_1149_));
 sg13g2_buf_2 fanout35 (.A(net37),
    .X(net35));
 sg13g2_and3_1 _1902_ (.X(_0130_),
    .A(net97),
    .B(_1136_),
    .C(net52));
 sg13g2_inv_1 _1903_ (.Y(_1152_),
    .A(_0036_));
 sg13g2_nor4_1 _1904_ (.A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[8] ),
    .C(\simon1.tick_counter[10] ),
    .D(\simon1.tick_counter[11] ),
    .Y(_1153_));
 sg13g2_nor4_1 _1905_ (.A(\simon1.tick_counter[12] ),
    .B(\simon1.tick_counter[13] ),
    .C(\simon1.tick_counter[14] ),
    .D(\simon1.tick_counter[15] ),
    .Y(_1154_));
 sg13g2_nor4_1 _1906_ (.A(\simon1.tick_counter[2] ),
    .B(\simon1.tick_counter[3] ),
    .C(\simon1.tick_counter[6] ),
    .D(\simon1.tick_counter[7] ),
    .Y(_1155_));
 sg13g2_inv_1 _1907_ (.Y(_1156_),
    .A(\simon1.tick_counter[0] ));
 sg13g2_nand2_1 _1908_ (.Y(_1157_),
    .A(\simon1.tick_counter[4] ),
    .B(\simon1.tick_counter[5] ));
 sg13g2_nor3_1 _1909_ (.A(_1156_),
    .B(\simon1.tick_counter[9] ),
    .C(_1157_),
    .Y(_1158_));
 sg13g2_and4_1 _1910_ (.A(_1153_),
    .B(_1154_),
    .C(_1155_),
    .D(_1158_),
    .X(_1159_));
 sg13g2_buf_1 fanout34 (.A(_0941_),
    .X(net34));
 sg13g2_nand2b_1 _1912_ (.Y(_1161_),
    .B(net95),
    .A_N(_1159_));
 sg13g2_buf_2 fanout33 (.A(net34),
    .X(net33));
 sg13g2_buf_2 fanout32 (.A(net34),
    .X(net32));
 sg13g2_nor2_1 _1915_ (.A(_1152_),
    .B(net40),
    .Y(_0161_));
 sg13g2_xnor2_1 _1916_ (.Y(_1164_),
    .A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[0] ));
 sg13g2_nor2_1 _1917_ (.A(net40),
    .B(_1164_),
    .Y(_0162_));
 sg13g2_nand2_1 _1918_ (.Y(_1165_),
    .A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[0] ));
 sg13g2_xor2_1 _1919_ (.B(_1165_),
    .A(\simon1.tick_counter[2] ),
    .X(_1166_));
 sg13g2_nor2_1 _1920_ (.A(net40),
    .B(_1166_),
    .Y(_0163_));
 sg13g2_nand3_1 _1921_ (.B(\simon1.tick_counter[0] ),
    .C(\simon1.tick_counter[2] ),
    .A(\simon1.tick_counter[1] ),
    .Y(_1167_));
 sg13g2_xor2_1 _1922_ (.B(_1167_),
    .A(\simon1.tick_counter[3] ),
    .X(_1168_));
 sg13g2_nor2_1 _1923_ (.A(net40),
    .B(_1168_),
    .Y(_0164_));
 sg13g2_inv_1 _1924_ (.Y(_1169_),
    .A(\simon1.tick_counter[4] ));
 sg13g2_nand4_1 _1925_ (.B(\simon1.tick_counter[0] ),
    .C(\simon1.tick_counter[2] ),
    .A(\simon1.tick_counter[1] ),
    .Y(_1170_),
    .D(\simon1.tick_counter[3] ));
 sg13g2_xnor2_1 _1926_ (.Y(_1171_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_nor2_1 _1927_ (.A(net40),
    .B(_1171_),
    .Y(_0165_));
 sg13g2_nor2_1 _1928_ (.A(_1169_),
    .B(_1170_),
    .Y(_1172_));
 sg13g2_xnor2_1 _1929_ (.Y(_1173_),
    .A(\simon1.tick_counter[5] ),
    .B(_1172_));
 sg13g2_nor2_1 _1930_ (.A(net40),
    .B(_1173_),
    .Y(_0166_));
 sg13g2_nor2_1 _1931_ (.A(_1157_),
    .B(_1170_),
    .Y(_1174_));
 sg13g2_xnor2_1 _1932_ (.Y(_1175_),
    .A(\simon1.tick_counter[6] ),
    .B(_1174_));
 sg13g2_nor2_1 _1933_ (.A(net39),
    .B(_1175_),
    .Y(_0167_));
 sg13g2_nand2_1 _1934_ (.Y(_1176_),
    .A(\simon1.tick_counter[6] ),
    .B(_1174_));
 sg13g2_xor2_1 _1935_ (.B(_1176_),
    .A(\simon1.tick_counter[7] ),
    .X(_1177_));
 sg13g2_nor2_1 _1936_ (.A(net39),
    .B(_1177_),
    .Y(_0168_));
 sg13g2_inv_1 _1937_ (.Y(_1178_),
    .A(\simon1.tick_counter[8] ));
 sg13g2_nand3_1 _1938_ (.B(\simon1.tick_counter[7] ),
    .C(_1174_),
    .A(\simon1.tick_counter[6] ),
    .Y(_1179_));
 sg13g2_xnor2_1 _1939_ (.Y(_1180_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_nor2_1 _1940_ (.A(net39),
    .B(_1180_),
    .Y(_0169_));
 sg13g2_nor2_1 _1941_ (.A(_1178_),
    .B(_1179_),
    .Y(_1181_));
 sg13g2_xnor2_1 _1942_ (.Y(_1182_),
    .A(\simon1.tick_counter[9] ),
    .B(_1181_));
 sg13g2_nor2_1 _1943_ (.A(net40),
    .B(_1182_),
    .Y(_0170_));
 sg13g2_nand2_1 _1944_ (.Y(_1183_),
    .A(\simon1.tick_counter[9] ),
    .B(_1181_));
 sg13g2_xor2_1 _1945_ (.B(_1183_),
    .A(\simon1.tick_counter[10] ),
    .X(_1184_));
 sg13g2_nor2_1 _1946_ (.A(net39),
    .B(_1184_),
    .Y(_0171_));
 sg13g2_inv_1 _1947_ (.Y(_1185_),
    .A(\simon1.tick_counter[11] ));
 sg13g2_nand3_1 _1948_ (.B(\simon1.tick_counter[10] ),
    .C(_1181_),
    .A(\simon1.tick_counter[9] ),
    .Y(_1186_));
 sg13g2_xnor2_1 _1949_ (.Y(_1187_),
    .A(_1185_),
    .B(_1186_));
 sg13g2_nor2_1 _1950_ (.A(net39),
    .B(_1187_),
    .Y(_0172_));
 sg13g2_nor2_2 _1951_ (.A(_1185_),
    .B(_1186_),
    .Y(_1188_));
 sg13g2_xnor2_1 _1952_ (.Y(_1189_),
    .A(\simon1.tick_counter[12] ),
    .B(_1188_));
 sg13g2_nor2_1 _1953_ (.A(net39),
    .B(_1189_),
    .Y(_0173_));
 sg13g2_nand2_1 _1954_ (.Y(_1190_),
    .A(\simon1.tick_counter[12] ),
    .B(_1188_));
 sg13g2_xor2_1 _1955_ (.B(_1190_),
    .A(\simon1.tick_counter[13] ),
    .X(_1191_));
 sg13g2_nor2_1 _1956_ (.A(net39),
    .B(_1191_),
    .Y(_0174_));
 sg13g2_nand3_1 _1957_ (.B(\simon1.tick_counter[13] ),
    .C(_1188_),
    .A(\simon1.tick_counter[12] ),
    .Y(_1192_));
 sg13g2_xor2_1 _1958_ (.B(_1192_),
    .A(\simon1.tick_counter[14] ),
    .X(_1193_));
 sg13g2_nor2_1 _1959_ (.A(_1161_),
    .B(_1193_),
    .Y(_0175_));
 sg13g2_nand4_1 _1960_ (.B(\simon1.tick_counter[13] ),
    .C(\simon1.tick_counter[14] ),
    .A(\simon1.tick_counter[12] ),
    .Y(_1194_),
    .D(_1188_));
 sg13g2_xor2_1 _1961_ (.B(_1194_),
    .A(\simon1.tick_counter[15] ),
    .X(_1195_));
 sg13g2_nor2_1 _1962_ (.A(net39),
    .B(_1195_),
    .Y(_0176_));
 sg13g2_nor2_2 _1963_ (.A(_0833_),
    .B(net43),
    .Y(_1196_));
 sg13g2_nand2_1 _1964_ (.Y(_1197_),
    .A(_0908_),
    .B(_1196_));
 sg13g2_nor2_1 _1965_ (.A(_0835_),
    .B(_1196_),
    .Y(_1198_));
 sg13g2_nor4_1 _1966_ (.A(_0859_),
    .B(_0922_),
    .C(_0933_),
    .D(_1198_),
    .Y(_1199_));
 sg13g2_o21ai_1 _1967_ (.B1(_1199_),
    .Y(_1200_),
    .A1(_0031_),
    .A2(_1197_));
 sg13g2_buf_1 fanout31 (.A(net34),
    .X(net31));
 sg13g2_a21oi_1 _1969_ (.A1(\simon1.state[6] ),
    .A2(_0929_),
    .Y(_1202_),
    .B1(net62));
 sg13g2_or3_1 _1970_ (.A(\simon1.seq_counter[0] ),
    .B(_1200_),
    .C(_1202_),
    .X(_1203_));
 sg13g2_nand2_1 _1971_ (.Y(_1204_),
    .A(\simon1.seq_counter[0] ),
    .B(_1200_));
 sg13g2_a21oi_1 _1972_ (.A1(_1203_),
    .A2(_1204_),
    .Y(_0082_),
    .B1(net86));
 sg13g2_a21oi_1 _1973_ (.A1(_0031_),
    .A2(_0908_),
    .Y(_1205_),
    .B1(_0853_));
 sg13g2_nor2_1 _1974_ (.A(_0835_),
    .B(_0031_),
    .Y(_1206_));
 sg13g2_o21ai_1 _1975_ (.B1(net95),
    .Y(_1207_),
    .A1(_1205_),
    .A2(_1206_));
 sg13g2_or2_1 _1976_ (.X(_1208_),
    .B(_1207_),
    .A(_1200_));
 sg13g2_buf_1 fanout30 (.A(net34),
    .X(net30));
 sg13g2_and2_1 _1978_ (.A(net95),
    .B(_1200_),
    .X(_1210_));
 sg13g2_buf_1 fanout29 (.A(_0953_),
    .X(net29));
 sg13g2_nor2_1 _1980_ (.A(\simon1.seq_counter[0] ),
    .B(_1207_),
    .Y(_1212_));
 sg13g2_o21ai_1 _1981_ (.B1(\simon1.seq_counter[1] ),
    .Y(_1213_),
    .A1(_1210_),
    .A2(_1212_));
 sg13g2_o21ai_1 _1982_ (.B1(_1213_),
    .Y(_0083_),
    .A1(_0884_),
    .A2(_1208_));
 sg13g2_nand2b_1 _1983_ (.Y(_1214_),
    .B(_0891_),
    .A_N(\simon1.seq_counter[2] ));
 sg13g2_nor2_1 _1984_ (.A(_0891_),
    .B(_1207_),
    .Y(_1215_));
 sg13g2_o21ai_1 _1985_ (.B1(\simon1.seq_counter[2] ),
    .Y(_1216_),
    .A1(_1210_),
    .A2(_1215_));
 sg13g2_o21ai_1 _1986_ (.B1(_1216_),
    .Y(_0084_),
    .A1(_1208_),
    .A2(_1214_));
 sg13g2_nand2b_1 _1987_ (.Y(_1217_),
    .B(_0895_),
    .A_N(\simon1.seq_counter[3] ));
 sg13g2_nor2_1 _1988_ (.A(_0895_),
    .B(_1207_),
    .Y(_1218_));
 sg13g2_o21ai_1 _1989_ (.B1(\simon1.seq_counter[3] ),
    .Y(_1219_),
    .A1(_1210_),
    .A2(_1218_));
 sg13g2_o21ai_1 _1990_ (.B1(_1219_),
    .Y(_0085_),
    .A1(_1208_),
    .A2(_1217_));
 sg13g2_nand2b_1 _1991_ (.Y(_1220_),
    .B(_0902_),
    .A_N(\simon1.seq_counter[4] ));
 sg13g2_nor2_1 _1992_ (.A(_0902_),
    .B(_1207_),
    .Y(_1221_));
 sg13g2_o21ai_1 _1993_ (.B1(\simon1.seq_counter[4] ),
    .Y(_1222_),
    .A1(_1210_),
    .A2(_1221_));
 sg13g2_o21ai_1 _1994_ (.B1(_1222_),
    .Y(_0086_),
    .A1(_1208_),
    .A2(_1220_));
 sg13g2_xnor2_1 _1995_ (.Y(_1223_),
    .A(\simon1.play1.tick_counter[0] ),
    .B(\simon1.play1.freq[0] ));
 sg13g2_nor2_1 _1996_ (.A(net89),
    .B(_1223_),
    .Y(_0098_));
 sg13g2_nand2_1 _1997_ (.Y(_1224_),
    .A(\simon1.play1.tick_counter[0] ),
    .B(\simon1.play1.freq[0] ));
 sg13g2_xnor2_1 _1998_ (.Y(_1225_),
    .A(\simon1.play1.tick_counter[1] ),
    .B(\simon1.play1.freq[1] ));
 sg13g2_xnor2_1 _1999_ (.Y(_1226_),
    .A(_1224_),
    .B(_1225_));
 sg13g2_nor2_1 _2000_ (.A(net89),
    .B(_1226_),
    .Y(_0099_));
 sg13g2_nor2_2 _2001_ (.A(\simon1.play1.tick_counter[1] ),
    .B(\simon1.play1.freq[1] ),
    .Y(_1227_));
 sg13g2_a22oi_1 _2002_ (.Y(_1228_),
    .B1(\simon1.play1.tick_counter[1] ),
    .B2(\simon1.play1.freq[1] ),
    .A2(\simon1.play1.freq[0] ),
    .A1(\simon1.play1.tick_counter[0] ));
 sg13g2_nor2_1 _2003_ (.A(_1227_),
    .B(_1228_),
    .Y(_1229_));
 sg13g2_xnor2_1 _2004_ (.Y(_1230_),
    .A(\simon1.play1.tick_counter[2] ),
    .B(\simon1.play1.freq[2] ));
 sg13g2_xor2_1 _2005_ (.B(_1230_),
    .A(_1229_),
    .X(_1231_));
 sg13g2_nor2_1 _2006_ (.A(net89),
    .B(_1231_),
    .Y(_0100_));
 sg13g2_and4_1 _2007_ (.A(_1139_),
    .B(_1142_),
    .C(_1145_),
    .D(_1149_),
    .X(_1232_));
 sg13g2_buf_2 fanout28 (.A(net29),
    .X(net28));
 sg13g2_buf_2 fanout27 (.A(net29),
    .X(net27));
 sg13g2_inv_1 _2010_ (.Y(_0213_),
    .A(\simon1.play1.freq[2] ));
 sg13g2_o21ai_1 _2011_ (.B1(_0213_),
    .Y(_0214_),
    .A1(_1227_),
    .A2(_1228_));
 sg13g2_nor3_1 _2012_ (.A(_0213_),
    .B(_1227_),
    .C(_1228_),
    .Y(_0215_));
 sg13g2_a21oi_1 _2013_ (.A1(\simon1.play1.tick_counter[2] ),
    .A2(_0214_),
    .Y(_0216_),
    .B1(_0215_));
 sg13g2_xor2_1 _2014_ (.B(_0216_),
    .A(\simon1.play1.freq[3] ),
    .X(_0217_));
 sg13g2_xnor2_1 _2015_ (.Y(_0218_),
    .A(_1134_),
    .B(_0217_));
 sg13g2_nor2_1 _2016_ (.A(net48),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_xnor2_1 _2017_ (.Y(_0220_),
    .A(\simon1.play1.tick_counter[3] ),
    .B(_0219_));
 sg13g2_nor2_1 _2018_ (.A(net89),
    .B(_0220_),
    .Y(_0101_));
 sg13g2_inv_1 _2019_ (.Y(_0221_),
    .A(\simon1.play1.tick_counter[4] ));
 sg13g2_nand2_2 _2020_ (.Y(_0222_),
    .A(_1119_),
    .B(_1133_));
 sg13g2_inv_1 _2021_ (.Y(_0223_),
    .A(\simon1.play1.tick_counter[3] ));
 sg13g2_xnor2_1 _2022_ (.Y(_0224_),
    .A(_0223_),
    .B(_0217_));
 sg13g2_nand2_1 _2023_ (.Y(_0225_),
    .A(_0222_),
    .B(_0224_));
 sg13g2_xnor2_1 _2024_ (.Y(_0226_),
    .A(\simon1.play1.tick_counter[3] ),
    .B(\simon1.play1.freq[3] ));
 sg13g2_nor4_2 _2025_ (.A(_1227_),
    .B(_1228_),
    .C(_1230_),
    .Y(_0227_),
    .D(_0226_));
 sg13g2_a21o_1 _2026_ (.A2(\simon1.play1.freq[2] ),
    .A1(\simon1.play1.tick_counter[2] ),
    .B1(\simon1.play1.freq[3] ),
    .X(_0228_));
 sg13g2_and3_1 _2027_ (.X(_0229_),
    .A(\simon1.play1.tick_counter[2] ),
    .B(\simon1.play1.freq[3] ),
    .C(\simon1.play1.freq[2] ));
 sg13g2_a21o_1 _2028_ (.A2(_0228_),
    .A1(\simon1.play1.tick_counter[3] ),
    .B1(_0229_),
    .X(_0230_));
 sg13g2_nor3_1 _2029_ (.A(\simon1.play1.freq[4] ),
    .B(_0227_),
    .C(_0230_),
    .Y(_0231_));
 sg13g2_or4_2 _2030_ (.A(_1227_),
    .B(_1228_),
    .C(_1230_),
    .D(_0226_),
    .X(_0232_));
 sg13g2_buf_1 fanout26 (.A(net29),
    .X(net26));
 sg13g2_a21oi_2 _2032_ (.B1(_0229_),
    .Y(_0234_),
    .A2(_0228_),
    .A1(\simon1.play1.tick_counter[3] ));
 sg13g2_inv_1 _2033_ (.Y(_0235_),
    .A(\simon1.play1.freq[4] ));
 sg13g2_a21oi_1 _2034_ (.A1(_0232_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_nor2_1 _2035_ (.A(_0231_),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_xnor2_1 _2036_ (.Y(_0238_),
    .A(_0225_),
    .B(_0237_));
 sg13g2_nand2_1 _2037_ (.Y(_0239_),
    .A(net52),
    .B(_0238_));
 sg13g2_xnor2_1 _2038_ (.Y(_0240_),
    .A(_0221_),
    .B(_0239_));
 sg13g2_nor2_1 _2039_ (.A(net91),
    .B(_0240_),
    .Y(_0102_));
 sg13g2_buf_1 fanout25 (.A(net29),
    .X(net25));
 sg13g2_buf_2 fanout24 (.A(_0462_),
    .X(net24));
 sg13g2_xor2_1 _2042_ (.B(net81),
    .A(net73),
    .X(_0243_));
 sg13g2_and2_1 _2043_ (.A(\simon1.play1.tick_counter[3] ),
    .B(_0228_),
    .X(_0244_));
 sg13g2_nor4_1 _2044_ (.A(\simon1.play1.tick_counter[4] ),
    .B(_0227_),
    .C(_0229_),
    .D(_0244_),
    .Y(_0245_));
 sg13g2_nor2_1 _2045_ (.A(\simon1.play1.tick_counter[4] ),
    .B(\simon1.play1.freq[4] ),
    .Y(_0246_));
 sg13g2_nor4_1 _2046_ (.A(_0231_),
    .B(_0243_),
    .C(_0245_),
    .D(_0246_),
    .Y(_0247_));
 sg13g2_nand3_1 _2047_ (.B(_0232_),
    .C(_0234_),
    .A(_0235_),
    .Y(_0248_));
 sg13g2_nand2b_1 _2048_ (.Y(_0249_),
    .B(net73),
    .A_N(net81));
 sg13g2_nand2b_1 _2049_ (.Y(_0250_),
    .B(net81),
    .A_N(net73));
 sg13g2_a221oi_1 _2050_ (.B2(_0250_),
    .C1(_0236_),
    .B1(_0249_),
    .A1(\simon1.play1.tick_counter[4] ),
    .Y(_0251_),
    .A2(_0248_));
 sg13g2_nor2_1 _2051_ (.A(_0247_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_xor2_1 _2052_ (.B(\simon1.play1.freq[4] ),
    .A(\simon1.play1.tick_counter[4] ),
    .X(_0253_));
 sg13g2_nand2b_1 _2053_ (.Y(_0254_),
    .B(_0253_),
    .A_N(_0226_));
 sg13g2_and2_1 _2054_ (.A(\simon1.play1.tick_counter[3] ),
    .B(\simon1.play1.freq[3] ),
    .X(_0255_));
 sg13g2_nor2_1 _2055_ (.A(\simon1.play1.freq[3] ),
    .B(_0253_),
    .Y(_0256_));
 sg13g2_a22oi_1 _2056_ (.Y(_0257_),
    .B1(_0256_),
    .B2(_0223_),
    .A2(_0255_),
    .A1(_0253_));
 sg13g2_mux2_1 _2057_ (.A0(_0254_),
    .A1(_0257_),
    .S(_0216_),
    .X(_0258_));
 sg13g2_nand2_1 _2058_ (.Y(_0259_),
    .A(_0222_),
    .B(_0258_));
 sg13g2_xnor2_1 _2059_ (.Y(_0260_),
    .A(_0252_),
    .B(_0259_));
 sg13g2_nor2_1 _2060_ (.A(net50),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_a21oi_1 _2061_ (.A1(net73),
    .A2(net50),
    .Y(_0262_),
    .B1(_0261_));
 sg13g2_nor2_1 _2062_ (.A(net91),
    .B(_0262_),
    .Y(_0103_));
 sg13g2_buf_2 fanout23 (.A(_0679_),
    .X(net23));
 sg13g2_o21ai_1 _2064_ (.B1(_0258_),
    .Y(_0264_),
    .A1(_0247_),
    .A2(_0251_));
 sg13g2_nand2_1 _2065_ (.Y(_0265_),
    .A(_0222_),
    .B(_0264_));
 sg13g2_nor2_1 _2066_ (.A(\simon1.play1.tick_counter[5] ),
    .B(\simon1.play1.freq[5] ),
    .Y(_0266_));
 sg13g2_a22oi_1 _2067_ (.Y(_0267_),
    .B1(\simon1.play1.freq[4] ),
    .B2(\simon1.play1.tick_counter[4] ),
    .A2(net81),
    .A1(\simon1.play1.tick_counter[5] ));
 sg13g2_nor2_2 _2068_ (.A(_0266_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_xnor2_1 _2069_ (.Y(_0269_),
    .A(\simon1.play1.tick_counter[4] ),
    .B(\simon1.play1.freq[4] ));
 sg13g2_a221oi_1 _2070_ (.B2(_0250_),
    .C1(_0269_),
    .B1(_0249_),
    .A1(_0232_),
    .Y(_0270_),
    .A2(_0234_));
 sg13g2_nor2_2 _2071_ (.A(_0268_),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_xor2_1 _2072_ (.B(_0271_),
    .A(net79),
    .X(_0272_));
 sg13g2_xnor2_1 _2073_ (.Y(_0273_),
    .A(_0265_),
    .B(_0272_));
 sg13g2_nor2_1 _2074_ (.A(net50),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_xnor2_1 _2075_ (.Y(_0275_),
    .A(\simon1.play1.tick_counter[6] ),
    .B(_0274_));
 sg13g2_nor2_1 _2076_ (.A(net92),
    .B(_0275_),
    .Y(_0104_));
 sg13g2_nor2_1 _2077_ (.A(\simon1.play1.tick_counter[7] ),
    .B(_1150_),
    .Y(_0276_));
 sg13g2_nand3_1 _2078_ (.B(_0232_),
    .C(_0234_),
    .A(\simon1.play1.freq[4] ),
    .Y(_0277_));
 sg13g2_xor2_1 _2079_ (.B(\simon1.play1.freq[7] ),
    .A(\simon1.play1.tick_counter[7] ),
    .X(_0278_));
 sg13g2_xor2_1 _2080_ (.B(net79),
    .A(\simon1.play1.tick_counter[6] ),
    .X(_0279_));
 sg13g2_nand3_1 _2081_ (.B(_0278_),
    .C(_0279_),
    .A(_0243_),
    .Y(_0280_));
 sg13g2_o21ai_1 _2082_ (.B1(_0280_),
    .Y(_0281_),
    .A1(_0227_),
    .A2(_0230_));
 sg13g2_a21oi_1 _2083_ (.A1(_0277_),
    .A2(_0281_),
    .Y(_0282_),
    .B1(_0221_));
 sg13g2_and2_1 _2084_ (.A(net73),
    .B(\simon1.play1.freq[5] ),
    .X(_0283_));
 sg13g2_a21oi_1 _2085_ (.A1(net79),
    .A2(_0283_),
    .Y(_0284_),
    .B1(\simon1.play1.tick_counter[6] ));
 sg13g2_nor2_1 _2086_ (.A(net79),
    .B(_0283_),
    .Y(_0285_));
 sg13g2_xnor2_1 _2087_ (.Y(_0286_),
    .A(\simon1.play1.tick_counter[7] ),
    .B(\simon1.play1.freq[7] ));
 sg13g2_o21ai_1 _2088_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_a21o_1 _2089_ (.A2(_0234_),
    .A1(_0232_),
    .B1(_0246_),
    .X(_0288_));
 sg13g2_xnor2_1 _2090_ (.Y(_0289_),
    .A(\simon1.play1.tick_counter[6] ),
    .B(net80));
 sg13g2_nor2_1 _2091_ (.A(_0286_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_a221oi_1 _2092_ (.B2(_0290_),
    .C1(_0235_),
    .B1(_0243_),
    .A1(_0232_),
    .Y(_0291_),
    .A2(_0234_));
 sg13g2_a21o_1 _2093_ (.A2(_0288_),
    .A1(_0287_),
    .B1(_0291_),
    .X(_0292_));
 sg13g2_o21ai_1 _2094_ (.B1(\simon1.play1.tick_counter[6] ),
    .Y(_0293_),
    .A1(net80),
    .A2(_0268_));
 sg13g2_a21oi_1 _2095_ (.A1(net79),
    .A2(_0268_),
    .Y(_0294_),
    .B1(_0286_));
 sg13g2_nor3_1 _2096_ (.A(net73),
    .B(net81),
    .C(net79),
    .Y(_0295_));
 sg13g2_o21ai_1 _2097_ (.B1(net79),
    .Y(_0296_),
    .A1(net73),
    .A2(net81));
 sg13g2_nor2b_1 _2098_ (.A(\simon1.play1.tick_counter[6] ),
    .B_N(_0296_),
    .Y(_0297_));
 sg13g2_nor3_1 _2099_ (.A(_0278_),
    .B(_0295_),
    .C(_0297_),
    .Y(_0298_));
 sg13g2_a21o_1 _2100_ (.A2(_0294_),
    .A1(_0293_),
    .B1(_0298_),
    .X(_0299_));
 sg13g2_o21ai_1 _2101_ (.B1(_0299_),
    .Y(_0300_),
    .A1(_0282_),
    .A2(_0292_));
 sg13g2_xnor2_1 _2102_ (.Y(_0301_),
    .A(_0271_),
    .B(_0289_));
 sg13g2_nand2_1 _2103_ (.Y(_0302_),
    .A(_0264_),
    .B(_0301_));
 sg13g2_and2_1 _2104_ (.A(_0222_),
    .B(_0302_),
    .X(_0303_));
 sg13g2_xnor2_1 _2105_ (.Y(_0304_),
    .A(_0300_),
    .B(_0303_));
 sg13g2_nor2_1 _2106_ (.A(net51),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_nor3_1 _2107_ (.A(net92),
    .B(_0276_),
    .C(_0305_),
    .Y(_0105_));
 sg13g2_nand4_1 _2108_ (.B(_0253_),
    .C(_0278_),
    .A(_0243_),
    .Y(_0306_),
    .D(_0279_));
 sg13g2_a21oi_2 _2109_ (.B1(_0306_),
    .Y(_0307_),
    .A2(_0234_),
    .A1(_0232_));
 sg13g2_nor2_1 _2110_ (.A(\simon1.play1.tick_counter[7] ),
    .B(\simon1.play1.freq[7] ),
    .Y(_0308_));
 sg13g2_a22oi_1 _2111_ (.Y(_0309_),
    .B1(net79),
    .B2(\simon1.play1.tick_counter[6] ),
    .A2(\simon1.play1.freq[7] ),
    .A1(\simon1.play1.tick_counter[7] ));
 sg13g2_or2_1 _2112_ (.X(_0310_),
    .B(_0309_),
    .A(_0308_));
 sg13g2_buf_2 fanout22 (.A(_0592_),
    .X(net22));
 sg13g2_or4_1 _2114_ (.A(_0266_),
    .B(_0267_),
    .C(_0286_),
    .D(_0289_),
    .X(_0312_));
 sg13g2_buf_2 fanout21 (.A(_0592_),
    .X(net21));
 sg13g2_nand2_1 _2116_ (.Y(_0314_),
    .A(_0310_),
    .B(_0312_));
 sg13g2_o21ai_1 _2117_ (.B1(net77),
    .Y(_0315_),
    .A1(_0307_),
    .A2(_0314_));
 sg13g2_or3_1 _2118_ (.A(net77),
    .B(_0307_),
    .C(_0314_),
    .X(_0316_));
 sg13g2_and2_1 _2119_ (.A(_0315_),
    .B(_0316_),
    .X(_0317_));
 sg13g2_nor2_1 _2120_ (.A(_0282_),
    .B(_0292_),
    .Y(_0318_));
 sg13g2_nor2b_1 _2121_ (.A(_0318_),
    .B_N(_0299_),
    .Y(_0319_));
 sg13g2_nand2_1 _2122_ (.Y(_0320_),
    .A(_0319_),
    .B(_0303_));
 sg13g2_xor2_1 _2123_ (.B(_0320_),
    .A(_0317_),
    .X(_0321_));
 sg13g2_nor2_1 _2124_ (.A(net50),
    .B(_0321_),
    .Y(_0322_));
 sg13g2_xnor2_1 _2125_ (.Y(_0323_),
    .A(net72),
    .B(_0322_));
 sg13g2_nor2_1 _2126_ (.A(net92),
    .B(_0323_),
    .Y(_0106_));
 sg13g2_inv_1 _2127_ (.Y(_0324_),
    .A(net72));
 sg13g2_a21o_1 _2128_ (.A2(_0316_),
    .A1(_0315_),
    .B1(_0324_),
    .X(_0325_));
 sg13g2_nand3_1 _2129_ (.B(_0315_),
    .C(_0316_),
    .A(_0324_),
    .Y(_0326_));
 sg13g2_a221oi_1 _2130_ (.B2(_0326_),
    .C1(_0300_),
    .B1(_0325_),
    .A1(_0264_),
    .Y(_0327_),
    .A2(_0301_));
 sg13g2_xnor2_1 _2131_ (.Y(_0328_),
    .A(\simon1.play1.tick_counter[9] ),
    .B(\simon1.play1.freq[9] ));
 sg13g2_inv_1 _2132_ (.Y(_0329_),
    .A(net78));
 sg13g2_nor2_1 _2133_ (.A(_0307_),
    .B(_0314_),
    .Y(_0330_));
 sg13g2_nor2_1 _2134_ (.A(_0308_),
    .B(_0309_),
    .Y(_0331_));
 sg13g2_nor2_1 _2135_ (.A(net72),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_o21ai_1 _2136_ (.B1(net77),
    .Y(_0333_),
    .A1(_0290_),
    .A2(_0331_));
 sg13g2_and2_1 _2137_ (.A(_0324_),
    .B(_0333_),
    .X(_0334_));
 sg13g2_a221oi_1 _2138_ (.B2(_0271_),
    .C1(_0334_),
    .B1(_0332_),
    .A1(_0329_),
    .Y(_0335_),
    .A2(_0330_));
 sg13g2_xnor2_1 _2139_ (.Y(_0336_),
    .A(_0328_),
    .B(_0335_));
 sg13g2_o21ai_1 _2140_ (.B1(_0336_),
    .Y(_0337_),
    .A1(_1134_),
    .A2(_0327_));
 sg13g2_a21oi_1 _2141_ (.A1(_0325_),
    .A2(_0326_),
    .Y(_0338_),
    .B1(_0300_));
 sg13g2_nand2_1 _2142_ (.Y(_0339_),
    .A(_0302_),
    .B(_0338_));
 sg13g2_nor2_1 _2143_ (.A(_1134_),
    .B(_0336_),
    .Y(_0340_));
 sg13g2_nand2_1 _2144_ (.Y(_0341_),
    .A(_0339_),
    .B(_0340_));
 sg13g2_nand3_1 _2145_ (.B(_0337_),
    .C(_0341_),
    .A(_1150_),
    .Y(_0342_));
 sg13g2_inv_1 _2146_ (.Y(_0343_),
    .A(\simon1.play1.tick_counter[9] ));
 sg13g2_a21oi_1 _2147_ (.A1(_0343_),
    .A2(net51),
    .Y(_0344_),
    .B1(net92));
 sg13g2_and2_1 _2148_ (.A(_0342_),
    .B(_0344_),
    .X(_0107_));
 sg13g2_nand2_1 _2149_ (.Y(_0345_),
    .A(\simon1.play1.tick_counter[10] ),
    .B(net50));
 sg13g2_inv_1 _2150_ (.Y(_0346_),
    .A(\simon1.play1.freq[9] ));
 sg13g2_nor2_1 _2151_ (.A(net72),
    .B(net77),
    .Y(_0347_));
 sg13g2_nor4_1 _2152_ (.A(_0346_),
    .B(_0308_),
    .C(_0309_),
    .D(_0347_),
    .Y(_0348_));
 sg13g2_and3_1 _2153_ (.X(_0349_),
    .A(net72),
    .B(\simon1.play1.freq[9] ),
    .C(net77));
 sg13g2_or3_1 _2154_ (.A(\simon1.play1.tick_counter[9] ),
    .B(_0348_),
    .C(_0349_),
    .X(_0350_));
 sg13g2_a21oi_1 _2155_ (.A1(net72),
    .A2(net77),
    .Y(_0351_),
    .B1(\simon1.play1.freq[9] ));
 sg13g2_o21ai_1 _2156_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0310_),
    .A2(_0347_));
 sg13g2_xor2_1 _2157_ (.B(net77),
    .A(\simon1.play1.tick_counter[8] ),
    .X(_0353_));
 sg13g2_nand2b_1 _2158_ (.Y(_0354_),
    .B(_0353_),
    .A_N(_0328_));
 sg13g2_nor2_1 _2159_ (.A(_0280_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_a21oi_1 _2160_ (.A1(_0232_),
    .A2(_0234_),
    .Y(_0356_),
    .B1(_0269_));
 sg13g2_nor2_1 _2161_ (.A(_0312_),
    .B(_0354_),
    .Y(_0357_));
 sg13g2_a221oi_1 _2162_ (.B2(_0356_),
    .C1(_0357_),
    .B1(_0355_),
    .A1(_0350_),
    .Y(_0358_),
    .A2(_0352_));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[6]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[4]));
 sg13g2_xor2_1 _2166_ (.B(_0358_),
    .A(_0035_),
    .X(_0362_));
 sg13g2_xnor2_1 _2167_ (.Y(_0363_),
    .A(_0341_),
    .B(_0362_));
 sg13g2_nand2_1 _2168_ (.Y(_0364_),
    .A(net52),
    .B(_0363_));
 sg13g2_a21oi_1 _2169_ (.A1(_0345_),
    .A2(_0364_),
    .Y(_0108_),
    .B1(net92));
 sg13g2_nand4_1 _2170_ (.B(_0339_),
    .C(_0340_),
    .A(_0035_),
    .Y(_0365_),
    .D(net38));
 sg13g2_nor2_1 _2171_ (.A(_0035_),
    .B(net38),
    .Y(_0366_));
 sg13g2_nand2_1 _2172_ (.Y(_0367_),
    .A(_0341_),
    .B(_0366_));
 sg13g2_a21oi_1 _2173_ (.A1(_0365_),
    .A2(_0367_),
    .Y(_0368_),
    .B1(net50));
 sg13g2_xnor2_1 _2174_ (.Y(_0369_),
    .A(net76),
    .B(_0368_));
 sg13g2_nor2_1 _2175_ (.A(net92),
    .B(_0369_),
    .Y(_0109_));
 sg13g2_nand2_1 _2176_ (.Y(_0370_),
    .A(\simon1.play1.tick_counter[12] ),
    .B(net51));
 sg13g2_a21o_1 _2177_ (.A2(net77),
    .A1(net72),
    .B1(\simon1.play1.freq[9] ),
    .X(_0371_));
 sg13g2_a21oi_1 _2178_ (.A1(\simon1.play1.tick_counter[9] ),
    .A2(_0371_),
    .Y(_0372_),
    .B1(_0349_));
 sg13g2_nand3_1 _2179_ (.B(_0310_),
    .C(_0372_),
    .A(net75),
    .Y(_0373_));
 sg13g2_nor3_1 _2180_ (.A(_0268_),
    .B(_0270_),
    .C(_0373_),
    .Y(_0374_));
 sg13g2_nand3_1 _2181_ (.B(_0312_),
    .C(_0372_),
    .A(_0310_),
    .Y(_0375_));
 sg13g2_o21ai_1 _2182_ (.B1(\simon1.play1.freq[9] ),
    .Y(_0376_),
    .A1(\simon1.play1.tick_counter[8] ),
    .A2(net78));
 sg13g2_nor3_1 _2183_ (.A(\simon1.play1.tick_counter[8] ),
    .B(\simon1.play1.freq[9] ),
    .C(net78),
    .Y(_0377_));
 sg13g2_a21o_1 _2184_ (.A2(_0376_),
    .A1(_0343_),
    .B1(_0377_),
    .X(_0378_));
 sg13g2_nand2_1 _2185_ (.Y(_0379_),
    .A(net76),
    .B(\simon1.play1.tick_counter[10] ));
 sg13g2_nor3_1 _2186_ (.A(net75),
    .B(_0378_),
    .C(_0379_),
    .Y(_0380_));
 sg13g2_o21ai_1 _2187_ (.B1(_0380_),
    .Y(_0381_),
    .A1(_0307_),
    .A2(_0375_));
 sg13g2_or2_1 _2188_ (.X(_0382_),
    .B(_0379_),
    .A(_0378_));
 sg13g2_nor2_1 _2189_ (.A(_0343_),
    .B(_0351_),
    .Y(_0383_));
 sg13g2_nor4_1 _2190_ (.A(_0290_),
    .B(_0331_),
    .C(_0349_),
    .D(_0383_),
    .Y(_0384_));
 sg13g2_o21ai_1 _2191_ (.B1(net75),
    .Y(_0385_),
    .A1(_0382_),
    .A2(_0384_));
 sg13g2_nand3b_1 _2192_ (.B(_0381_),
    .C(_0385_),
    .Y(_0386_),
    .A_N(_0374_));
 sg13g2_nor2b_1 _2193_ (.A(_0035_),
    .B_N(\simon1.play1.tick_counter[11] ),
    .Y(_0387_));
 sg13g2_nor2b_1 _2194_ (.A(net76),
    .B_N(_0035_),
    .Y(_0388_));
 sg13g2_mux2_1 _2195_ (.A0(_0387_),
    .A1(_0388_),
    .S(net38),
    .X(_0389_));
 sg13g2_nand3_1 _2196_ (.B(_0340_),
    .C(_0389_),
    .A(_0339_),
    .Y(_0390_));
 sg13g2_xnor2_1 _2197_ (.Y(_0391_),
    .A(_0386_),
    .B(_0390_));
 sg13g2_nand2_1 _2198_ (.Y(_0392_),
    .A(_1150_),
    .B(_0391_));
 sg13g2_a21oi_1 _2199_ (.A1(_0370_),
    .A2(_0392_),
    .Y(_0110_),
    .B1(net92));
 sg13g2_nand2b_1 _2200_ (.Y(_0393_),
    .B(_0389_),
    .A_N(_0386_));
 sg13g2_or3_1 _2201_ (.A(_0336_),
    .B(_0327_),
    .C(_0393_),
    .X(_0394_));
 sg13g2_nand2_1 _2202_ (.Y(_0395_),
    .A(_0222_),
    .B(_0394_));
 sg13g2_nand2_2 _2203_ (.Y(_0396_),
    .A(net75),
    .B(_0387_));
 sg13g2_nor2_2 _2204_ (.A(net38),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_xor2_1 _2205_ (.B(_0397_),
    .A(_0395_),
    .X(_0398_));
 sg13g2_nor2_1 _2206_ (.A(net51),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_xnor2_1 _2207_ (.Y(_0400_),
    .A(\simon1.play1.tick_counter[13] ),
    .B(_0399_));
 sg13g2_nor2_1 _2208_ (.A(net93),
    .B(_0400_),
    .Y(_0111_));
 sg13g2_nand4_1 _2209_ (.B(\simon1.play1.tick_counter[13] ),
    .C(net76),
    .A(net75),
    .Y(_0401_),
    .D(\simon1.play1.tick_counter[10] ));
 sg13g2_nand2_1 _2210_ (.Y(_0402_),
    .A(_0396_),
    .B(_0401_));
 sg13g2_nand3b_1 _2211_ (.B(_0402_),
    .C(\simon1.play1.tick_counter[13] ),
    .Y(_0403_),
    .A_N(net38));
 sg13g2_o21ai_1 _2212_ (.B1(_0403_),
    .Y(_0404_),
    .A1(\simon1.play1.tick_counter[13] ),
    .A2(_0397_));
 sg13g2_or2_1 _2213_ (.X(_0405_),
    .B(_0404_),
    .A(_0395_));
 sg13g2_and2_1 _2214_ (.A(net75),
    .B(_0387_),
    .X(_0406_));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[3]));
 sg13g2_nor2_1 _2216_ (.A(net38),
    .B(_0401_),
    .Y(_0408_));
 sg13g2_o21ai_1 _2217_ (.B1(_0408_),
    .Y(_0409_),
    .A1(_0395_),
    .A2(_0406_));
 sg13g2_a21oi_1 _2218_ (.A1(_0405_),
    .A2(_0409_),
    .Y(_0410_),
    .B1(net50));
 sg13g2_xnor2_1 _2219_ (.Y(_0411_),
    .A(\simon1.play1.tick_counter[14] ),
    .B(_0410_));
 sg13g2_nor2_1 _2220_ (.A(net91),
    .B(_0411_),
    .Y(_0112_));
 sg13g2_nor2_1 _2221_ (.A(\simon1.play1.tick_counter[13] ),
    .B(_0397_),
    .Y(_0412_));
 sg13g2_nand2_1 _2222_ (.Y(_0413_),
    .A(\simon1.play1.tick_counter[14] ),
    .B(_0403_));
 sg13g2_nand3b_1 _2223_ (.B(_0396_),
    .C(_0408_),
    .Y(_0414_),
    .A_N(\simon1.play1.tick_counter[14] ));
 sg13g2_o21ai_1 _2224_ (.B1(_0414_),
    .Y(_0415_),
    .A1(_0412_),
    .A2(_0413_));
 sg13g2_a21oi_2 _2225_ (.B1(_1134_),
    .Y(_0416_),
    .A2(_0415_),
    .A1(_0394_));
 sg13g2_a21oi_1 _2226_ (.A1(_1102_),
    .A2(_0397_),
    .Y(_0417_),
    .B1(net50));
 sg13g2_nand2_1 _2227_ (.Y(_0418_),
    .A(_0416_),
    .B(_0417_));
 sg13g2_xor2_1 _2228_ (.B(_0418_),
    .A(\simon1.play1.tick_counter[15] ),
    .X(_0419_));
 sg13g2_nor2_1 _2229_ (.A(net93),
    .B(_0419_),
    .Y(_0113_));
 sg13g2_nand2_1 _2230_ (.Y(_0420_),
    .A(\simon1.play1.tick_counter[16] ),
    .B(net48));
 sg13g2_nand3_1 _2231_ (.B(\simon1.play1.tick_counter[10] ),
    .C(_0349_),
    .A(net76),
    .Y(_0421_));
 sg13g2_nand4_1 _2232_ (.B(\simon1.play1.tick_counter[10] ),
    .C(\simon1.play1.tick_counter[9] ),
    .A(net76),
    .Y(_0422_),
    .D(_0371_));
 sg13g2_nand4_1 _2233_ (.B(_0312_),
    .C(_0421_),
    .A(_0310_),
    .Y(_0423_),
    .D(_0422_));
 sg13g2_and3_1 _2234_ (.X(_0424_),
    .A(net75),
    .B(net76),
    .C(\simon1.play1.tick_counter[10] ));
 sg13g2_nand3_1 _2235_ (.B(_1102_),
    .C(_0424_),
    .A(\simon1.play1.tick_counter[15] ),
    .Y(_0425_));
 sg13g2_nor2_1 _2236_ (.A(_0378_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_o21ai_1 _2237_ (.B1(_0426_),
    .Y(_0427_),
    .A1(_0307_),
    .A2(_0423_));
 sg13g2_xor2_1 _2238_ (.B(_0427_),
    .A(\simon1.play1.tick_counter[16] ),
    .X(_0428_));
 sg13g2_nand2_1 _2239_ (.Y(_0429_),
    .A(_1102_),
    .B(_0406_));
 sg13g2_o21ai_1 _2240_ (.B1(\simon1.play1.tick_counter[15] ),
    .Y(_0430_),
    .A1(net38),
    .A2(_0429_));
 sg13g2_or3_1 _2241_ (.A(\simon1.play1.tick_counter[15] ),
    .B(net38),
    .C(_0429_),
    .X(_0431_));
 sg13g2_nand3_1 _2242_ (.B(_0430_),
    .C(_0431_),
    .A(_0416_),
    .Y(_0432_));
 sg13g2_xor2_1 _2243_ (.B(_0432_),
    .A(_0428_),
    .X(_0433_));
 sg13g2_nand2_1 _2244_ (.Y(_0434_),
    .A(net52),
    .B(_0433_));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_a21oi_1 _2246_ (.A1(_0420_),
    .A2(_0434_),
    .Y(_0114_),
    .B1(net90));
 sg13g2_nand3_1 _2247_ (.B(\simon1.play1.tick_counter[16] ),
    .C(_1102_),
    .A(\simon1.play1.tick_counter[15] ),
    .Y(_0436_));
 sg13g2_or2_2 _2248_ (.X(_0437_),
    .B(_0436_),
    .A(_0396_));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_nor2_1 _2250_ (.A(net35),
    .B(_0437_),
    .Y(_0439_));
 sg13g2_nand4_1 _2251_ (.B(\simon1.play1.tick_counter[16] ),
    .C(_1102_),
    .A(\simon1.play1.tick_counter[15] ),
    .Y(_0440_),
    .D(_0424_));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_or2_1 _2253_ (.X(_0442_),
    .B(_0440_),
    .A(net37));
 sg13g2_nand2_1 _2254_ (.Y(_0443_),
    .A(_0439_),
    .B(_0442_));
 sg13g2_and3_1 _2255_ (.X(_0444_),
    .A(_0428_),
    .B(_0430_),
    .C(_0431_));
 sg13g2_or2_2 _2256_ (.X(_0445_),
    .B(_0437_),
    .A(net37));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_nand3_1 _2258_ (.B(_0444_),
    .C(_0445_),
    .A(_0416_),
    .Y(_0447_));
 sg13g2_a21oi_1 _2259_ (.A1(_0443_),
    .A2(_0447_),
    .Y(_0448_),
    .B1(net48));
 sg13g2_xnor2_1 _2260_ (.Y(_0449_),
    .A(\simon1.play1.tick_counter[17] ),
    .B(_0448_));
 sg13g2_nor2_1 _2261_ (.A(net90),
    .B(_0449_),
    .Y(_0115_));
 sg13g2_a21oi_1 _2262_ (.A1(_0428_),
    .A2(_0439_),
    .Y(_0450_),
    .B1(_0442_));
 sg13g2_nand2_1 _2263_ (.Y(_0451_),
    .A(\simon1.play1.tick_counter[17] ),
    .B(_0450_));
 sg13g2_nor2_1 _2264_ (.A(\simon1.play1.tick_counter[17] ),
    .B(_0439_),
    .Y(_0452_));
 sg13g2_nand3_1 _2265_ (.B(_0444_),
    .C(_0452_),
    .A(_0416_),
    .Y(_0453_));
 sg13g2_a21oi_1 _2266_ (.A1(_0451_),
    .A2(_0453_),
    .Y(_0454_),
    .B1(net48));
 sg13g2_xnor2_1 _2267_ (.Y(_0455_),
    .A(\simon1.play1.tick_counter[18] ),
    .B(_0454_));
 sg13g2_nor2_1 _2268_ (.A(net89),
    .B(_0455_),
    .Y(_0116_));
 sg13g2_nand2_1 _2269_ (.Y(_0456_),
    .A(\simon1.play1.tick_counter[18] ),
    .B(\simon1.play1.tick_counter[17] ));
 sg13g2_nor2_1 _2270_ (.A(_0445_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor2_1 _2271_ (.A(\simon1.play1.tick_counter[18] ),
    .B(\simon1.play1.tick_counter[17] ),
    .Y(_0458_));
 sg13g2_nor4_1 _2272_ (.A(net37),
    .B(_0437_),
    .C(net45),
    .D(_0456_),
    .Y(_0459_));
 sg13g2_a21o_1 _2273_ (.A2(_0445_),
    .A1(_0458_),
    .B1(_0459_),
    .X(_0460_));
 sg13g2_nand3_1 _2274_ (.B(_0444_),
    .C(_0460_),
    .A(_0222_),
    .Y(_0461_));
 sg13g2_a21oi_1 _2275_ (.A1(_0394_),
    .A2(_0415_),
    .Y(_0462_),
    .B1(_0461_));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_xnor2_1 _2277_ (.Y(_0464_),
    .A(_0457_),
    .B(_0462_));
 sg13g2_nor2_1 _2278_ (.A(net49),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_xnor2_1 _2279_ (.Y(_0466_),
    .A(\simon1.play1.tick_counter[19] ),
    .B(_0465_));
 sg13g2_nor2_1 _2280_ (.A(net93),
    .B(_0466_),
    .Y(_0117_));
 sg13g2_nand2_1 _2281_ (.Y(_0467_),
    .A(\simon1.play1.tick_counter[20] ),
    .B(net48));
 sg13g2_inv_1 _2282_ (.Y(_0468_),
    .A(\simon1.play1.tick_counter[19] ));
 sg13g2_nor4_1 _2283_ (.A(_0468_),
    .B(_0378_),
    .C(net45),
    .D(_0456_),
    .Y(_0469_));
 sg13g2_o21ai_1 _2284_ (.B1(_0469_),
    .Y(_0470_),
    .A1(_0307_),
    .A2(_0423_));
 sg13g2_xor2_1 _2285_ (.B(_0470_),
    .A(\simon1.play1.tick_counter[20] ),
    .X(_0471_));
 sg13g2_xnor2_1 _2286_ (.Y(_0472_),
    .A(\simon1.play1.tick_counter[19] ),
    .B(_0457_));
 sg13g2_nand2_1 _2287_ (.Y(_0473_),
    .A(net24),
    .B(_0472_));
 sg13g2_nand2b_1 _2288_ (.Y(_0474_),
    .B(_0473_),
    .A_N(_0471_));
 sg13g2_nand3_1 _2289_ (.B(_0471_),
    .C(_0472_),
    .A(net24),
    .Y(_0475_));
 sg13g2_a21o_1 _2290_ (.A2(_0475_),
    .A1(_0474_),
    .B1(net48),
    .X(_0476_));
 sg13g2_a21oi_1 _2291_ (.A1(_0467_),
    .A2(_0476_),
    .Y(_0118_),
    .B1(net89));
 sg13g2_nand4_1 _2292_ (.B(\simon1.play1.tick_counter[19] ),
    .C(\simon1.play1.tick_counter[18] ),
    .A(\simon1.play1.tick_counter[20] ),
    .Y(_0477_),
    .D(\simon1.play1.tick_counter[17] ));
 sg13g2_nor2_1 _2293_ (.A(_0445_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_xor2_1 _2294_ (.B(_0478_),
    .A(_0475_),
    .X(_0479_));
 sg13g2_o21ai_1 _2295_ (.B1(\simon1.play1.tick_counter[21] ),
    .Y(_0480_),
    .A1(net48),
    .A2(_0479_));
 sg13g2_or3_1 _2296_ (.A(\simon1.play1.tick_counter[21] ),
    .B(net48),
    .C(_0479_),
    .X(_0481_));
 sg13g2_a21oi_1 _2297_ (.A1(_0480_),
    .A2(_0481_),
    .Y(_0119_),
    .B1(net89));
 sg13g2_and2_1 _2298_ (.A(net96),
    .B(\simon1.play1.tick_counter[22] ),
    .X(_0482_));
 sg13g2_nor2_1 _2299_ (.A(net88),
    .B(\simon1.play1.tick_counter[22] ),
    .Y(_0483_));
 sg13g2_nor2_1 _2300_ (.A(net35),
    .B(net45),
    .Y(_0484_));
 sg13g2_inv_1 _2301_ (.Y(_0485_),
    .A(\simon1.play1.tick_counter[21] ));
 sg13g2_nor2_1 _2302_ (.A(_0485_),
    .B(_0477_),
    .Y(_0486_));
 sg13g2_nand2_1 _2303_ (.Y(_0487_),
    .A(_0484_),
    .B(_0486_));
 sg13g2_xnor2_1 _2304_ (.Y(_0488_),
    .A(\simon1.play1.tick_counter[21] ),
    .B(_0478_));
 sg13g2_nand4_1 _2305_ (.B(_0471_),
    .C(_0472_),
    .A(net24),
    .Y(_0489_),
    .D(_0488_));
 sg13g2_xnor2_1 _2306_ (.Y(_0490_),
    .A(_0487_),
    .B(_0489_));
 sg13g2_nor2_1 _2307_ (.A(net47),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_mux2_1 _2308_ (.A0(_0482_),
    .A1(_0483_),
    .S(_0491_),
    .X(_0120_));
 sg13g2_nand2_1 _2309_ (.Y(_0492_),
    .A(\simon1.play1.tick_counter[22] ),
    .B(_0486_));
 sg13g2_nor2_1 _2310_ (.A(_0445_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nor2_1 _2311_ (.A(_0436_),
    .B(_0477_),
    .Y(_0494_));
 sg13g2_nand2_1 _2312_ (.Y(_0495_),
    .A(_0406_),
    .B(_0494_));
 sg13g2_nor2_1 _2313_ (.A(\simon1.play1.tick_counter[22] ),
    .B(\simon1.play1.tick_counter[21] ),
    .Y(_0496_));
 sg13g2_o21ai_1 _2314_ (.B1(_0496_),
    .Y(_0497_),
    .A1(net35),
    .A2(_0495_));
 sg13g2_nand4_1 _2315_ (.B(_0406_),
    .C(net45),
    .A(\simon1.play1.tick_counter[21] ),
    .Y(_0498_),
    .D(_0494_));
 sg13g2_or3_1 _2316_ (.A(\simon1.play1.tick_counter[22] ),
    .B(net35),
    .C(_0498_),
    .X(_0499_));
 sg13g2_nand2_1 _2317_ (.Y(_0500_),
    .A(\simon1.play1.tick_counter[22] ),
    .B(\simon1.play1.tick_counter[21] ));
 sg13g2_or4_1 _2318_ (.A(net36),
    .B(net45),
    .C(_0495_),
    .D(_0500_),
    .X(_0501_));
 sg13g2_nand3_1 _2319_ (.B(_0499_),
    .C(_0501_),
    .A(_0497_),
    .Y(_0502_));
 sg13g2_nand4_1 _2320_ (.B(_0471_),
    .C(_0472_),
    .A(net24),
    .Y(_0503_),
    .D(_0502_));
 sg13g2_xnor2_1 _2321_ (.Y(_0504_),
    .A(_0493_),
    .B(_0503_));
 sg13g2_nand2_1 _2322_ (.Y(_0505_),
    .A(net96),
    .B(\simon1.play1.tick_counter[23] ));
 sg13g2_a21oi_1 _2323_ (.A1(net52),
    .A2(_0504_),
    .Y(_0506_),
    .B1(_0505_));
 sg13g2_inv_1 _2324_ (.Y(_0507_),
    .A(\simon1.play1.tick_counter[23] ));
 sg13g2_nand4_1 _2325_ (.B(_0507_),
    .C(net52),
    .A(net96),
    .Y(_0508_),
    .D(_0504_));
 sg13g2_nand2b_1 _2326_ (.Y(_0121_),
    .B(_0508_),
    .A_N(_0506_));
 sg13g2_nand2_1 _2327_ (.Y(_0509_),
    .A(\simon1.play1.tick_counter[24] ),
    .B(net47));
 sg13g2_nor4_1 _2328_ (.A(_0507_),
    .B(net35),
    .C(net45),
    .D(_0492_),
    .Y(_0510_));
 sg13g2_xnor2_1 _2329_ (.Y(_0511_),
    .A(\simon1.play1.tick_counter[24] ),
    .B(_0510_));
 sg13g2_nor4_1 _2330_ (.A(\simon1.play1.tick_counter[23] ),
    .B(net35),
    .C(_0437_),
    .D(_0492_),
    .Y(_0512_));
 sg13g2_o21ai_1 _2331_ (.B1(\simon1.play1.tick_counter[23] ),
    .Y(_0513_),
    .A1(_0445_),
    .A2(_0492_));
 sg13g2_nor2b_1 _2332_ (.A(_0512_),
    .B_N(_0513_),
    .Y(_0514_));
 sg13g2_and2_1 _2333_ (.A(_0502_),
    .B(_0514_),
    .X(_0515_));
 sg13g2_nand4_1 _2334_ (.B(_0471_),
    .C(_0472_),
    .A(net24),
    .Y(_0516_),
    .D(_0515_));
 sg13g2_xor2_1 _2335_ (.B(_0516_),
    .A(_0511_),
    .X(_0517_));
 sg13g2_nand2_1 _2336_ (.Y(_0518_),
    .A(net52),
    .B(_0517_));
 sg13g2_a21oi_1 _2337_ (.A1(_0509_),
    .A2(_0518_),
    .Y(_0122_),
    .B1(net88));
 sg13g2_nor2b_1 _2338_ (.A(_0512_),
    .B_N(_0471_),
    .Y(_0519_));
 sg13g2_nand4_1 _2339_ (.B(_0511_),
    .C(_0513_),
    .A(_0502_),
    .Y(_0520_),
    .D(_0519_));
 sg13g2_inv_1 _2340_ (.Y(_0521_),
    .A(_0520_));
 sg13g2_nand3_1 _2341_ (.B(_0472_),
    .C(_0521_),
    .A(net24),
    .Y(_0522_));
 sg13g2_nand4_1 _2342_ (.B(\simon1.play1.tick_counter[23] ),
    .C(\simon1.play1.tick_counter[22] ),
    .A(\simon1.play1.tick_counter[24] ),
    .Y(_0523_),
    .D(_0486_));
 sg13g2_nor3_2 _2343_ (.A(net35),
    .B(_0437_),
    .C(_0523_),
    .Y(_0524_));
 sg13g2_xor2_1 _2344_ (.B(_0524_),
    .A(_0522_),
    .X(_0525_));
 sg13g2_o21ai_1 _2345_ (.B1(\simon1.play1.tick_counter[25] ),
    .Y(_0526_),
    .A1(net46),
    .A2(_0525_));
 sg13g2_or3_1 _2346_ (.A(\simon1.play1.tick_counter[25] ),
    .B(net47),
    .C(_0525_),
    .X(_0527_));
 sg13g2_a21oi_1 _2347_ (.A1(_0526_),
    .A2(_0527_),
    .Y(_0123_),
    .B1(net88));
 sg13g2_nor2_1 _2348_ (.A(net88),
    .B(\simon1.play1.tick_counter[26] ),
    .Y(_0528_));
 sg13g2_inv_2 _2349_ (.Y(_0529_),
    .A(\simon1.play1.tick_counter[26] ));
 sg13g2_nor2_1 _2350_ (.A(net88),
    .B(_0529_),
    .Y(_0530_));
 sg13g2_inv_1 _2351_ (.Y(_0531_),
    .A(\simon1.play1.tick_counter[25] ));
 sg13g2_nor2_1 _2352_ (.A(_0531_),
    .B(net46),
    .Y(_0532_));
 sg13g2_nor4_1 _2353_ (.A(net35),
    .B(_0439_),
    .C(net45),
    .D(_0523_),
    .Y(_0533_));
 sg13g2_nor3_1 _2354_ (.A(\simon1.play1.tick_counter[25] ),
    .B(net47),
    .C(_0524_),
    .Y(_0534_));
 sg13g2_nor2_1 _2355_ (.A(_0473_),
    .B(_0520_),
    .Y(_0535_));
 sg13g2_a22oi_1 _2356_ (.Y(_0536_),
    .B1(_0534_),
    .B2(_0535_),
    .A2(_0533_),
    .A1(_0532_));
 sg13g2_mux2_1 _2357_ (.A0(_0528_),
    .A1(_0530_),
    .S(_0536_),
    .X(_0124_));
 sg13g2_nor2_1 _2358_ (.A(\simon1.play1.tick_counter[25] ),
    .B(_0524_),
    .Y(_0537_));
 sg13g2_nor4_1 _2359_ (.A(_0531_),
    .B(_0445_),
    .C(_0484_),
    .D(_0523_),
    .Y(_0538_));
 sg13g2_o21ai_1 _2360_ (.B1(_0529_),
    .Y(_0539_),
    .A1(_0537_),
    .A2(_0538_));
 sg13g2_and2_1 _2361_ (.A(\simon1.play1.tick_counter[25] ),
    .B(_0524_),
    .X(_0540_));
 sg13g2_nor2_1 _2362_ (.A(_0529_),
    .B(_0442_),
    .Y(_0541_));
 sg13g2_nand2_1 _2363_ (.Y(_0542_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_a21oi_1 _2364_ (.A1(_0539_),
    .A2(_0542_),
    .Y(_0543_),
    .B1(_0520_));
 sg13g2_nand3_1 _2365_ (.B(_0472_),
    .C(_0543_),
    .A(net24),
    .Y(_0544_));
 sg13g2_or2_1 _2366_ (.X(_0545_),
    .B(_0523_),
    .A(_0531_));
 sg13g2_nor4_2 _2367_ (.A(_0529_),
    .B(net36),
    .C(_0437_),
    .Y(_0546_),
    .D(_0545_));
 sg13g2_xor2_1 _2368_ (.B(_0546_),
    .A(_0544_),
    .X(_0547_));
 sg13g2_o21ai_1 _2369_ (.B1(net74),
    .Y(_0548_),
    .A1(net46),
    .A2(_0547_));
 sg13g2_or3_1 _2370_ (.A(net74),
    .B(net46),
    .C(_0547_),
    .X(_0549_));
 sg13g2_a21oi_1 _2371_ (.A1(_0548_),
    .A2(_0549_),
    .Y(_0125_),
    .B1(net88));
 sg13g2_inv_1 _2372_ (.Y(_0550_),
    .A(net74));
 sg13g2_nor4_2 _2373_ (.A(_0529_),
    .B(net36),
    .C(net45),
    .Y(_0551_),
    .D(_0545_));
 sg13g2_o21ai_1 _2374_ (.B1(net52),
    .Y(_0552_),
    .A1(_0550_),
    .A2(_0551_));
 sg13g2_a221oi_1 _2375_ (.B2(_0550_),
    .C1(_0552_),
    .B1(_0544_),
    .A1(_0540_),
    .Y(_0553_),
    .A2(_0541_));
 sg13g2_xnor2_1 _2376_ (.Y(_0554_),
    .A(\simon1.play1.tick_counter[28] ),
    .B(_0553_));
 sg13g2_nor2_1 _2377_ (.A(net88),
    .B(_0554_),
    .Y(_0126_));
 sg13g2_and2_1 _2378_ (.A(net96),
    .B(\simon1.play1.tick_counter[29] ),
    .X(_0555_));
 sg13g2_nor2_1 _2379_ (.A(net88),
    .B(\simon1.play1.tick_counter[29] ),
    .Y(_0556_));
 sg13g2_or4_1 _2380_ (.A(\simon1.play1.tick_counter[28] ),
    .B(net74),
    .C(_0544_),
    .D(_0546_),
    .X(_0557_));
 sg13g2_nand4_1 _2381_ (.B(net74),
    .C(_0544_),
    .A(\simon1.play1.tick_counter[28] ),
    .Y(_0558_),
    .D(_0546_));
 sg13g2_a21oi_1 _2382_ (.A1(_0557_),
    .A2(_0558_),
    .Y(_0559_),
    .B1(net46));
 sg13g2_mux2_1 _2383_ (.A0(_0555_),
    .A1(_0556_),
    .S(_0559_),
    .X(_0127_));
 sg13g2_and3_1 _2384_ (.X(_0560_),
    .A(\simon1.play1.tick_counter[29] ),
    .B(\simon1.play1.tick_counter[28] ),
    .C(\simon1.play1.tick_counter[27] ));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_nand2_1 _2386_ (.Y(_0562_),
    .A(_0551_),
    .B(_0560_));
 sg13g2_nor2b_1 _2387_ (.A(_0551_),
    .B_N(_0546_),
    .Y(_0563_));
 sg13g2_nor2_1 _2388_ (.A(net74),
    .B(_0546_),
    .Y(_0564_));
 sg13g2_a21oi_1 _2389_ (.A1(net74),
    .A2(_0563_),
    .Y(_0565_),
    .B1(_0564_));
 sg13g2_nand3_1 _2390_ (.B(_0551_),
    .C(_0560_),
    .A(_0546_),
    .Y(_0566_));
 sg13g2_o21ai_1 _2391_ (.B1(_0566_),
    .Y(_0567_),
    .A1(_1129_),
    .A2(_0565_));
 sg13g2_nand4_1 _2392_ (.B(_0472_),
    .C(_0543_),
    .A(net24),
    .Y(_0568_),
    .D(_0567_));
 sg13g2_xnor2_1 _2393_ (.Y(_0569_),
    .A(_0562_),
    .B(_0568_));
 sg13g2_o21ai_1 _2394_ (.B1(\simon1.play1.tick_counter[30] ),
    .Y(_0570_),
    .A1(net46),
    .A2(_0569_));
 sg13g2_or3_1 _2395_ (.A(\simon1.play1.tick_counter[30] ),
    .B(net46),
    .C(_0569_),
    .X(_0571_));
 sg13g2_a21oi_1 _2396_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0128_),
    .B1(net90));
 sg13g2_nand2_1 _2397_ (.Y(_0572_),
    .A(\simon1.play1.tick_counter[26] ),
    .B(_0406_));
 sg13g2_nor4_1 _2398_ (.A(net36),
    .B(_0436_),
    .C(_0545_),
    .D(_0572_),
    .Y(_0573_));
 sg13g2_nand3_1 _2399_ (.B(_0573_),
    .C(_0560_),
    .A(\simon1.play1.tick_counter[30] ),
    .Y(_0574_));
 sg13g2_o21ai_1 _2400_ (.B1(_0560_),
    .Y(_0575_),
    .A1(_0546_),
    .A2(_0551_));
 sg13g2_a21oi_1 _2401_ (.A1(\simon1.play1.tick_counter[30] ),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net46));
 sg13g2_nand2_1 _2402_ (.Y(_0577_),
    .A(_0566_),
    .B(_0576_));
 sg13g2_a21oi_1 _2403_ (.A1(_0568_),
    .A2(_0574_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_xnor2_1 _2404_ (.Y(_0579_),
    .A(\simon1.play1.tick_counter[31] ),
    .B(_0578_));
 sg13g2_nor2_1 _2405_ (.A(net90),
    .B(_0579_),
    .Y(_0129_));
 sg13g2_a21oi_1 _2406_ (.A1(\simon1.state[0] ),
    .A2(_0848_),
    .Y(_0580_),
    .B1(\simon1.score1.ena ));
 sg13g2_nor2_1 _2407_ (.A(net94),
    .B(_0580_),
    .Y(_0132_));
 sg13g2_nor3_1 _2408_ (.A(net86),
    .B(_0031_),
    .C(_1197_),
    .Y(_0133_));
 sg13g2_and2_1 _2409_ (.A(net95),
    .B(_0037_),
    .X(_0136_));
 sg13g2_xnor2_1 _2410_ (.Y(_0581_),
    .A(\simon1.next_random[1] ),
    .B(\simon1.next_random[0] ));
 sg13g2_nor2_1 _2411_ (.A(net87),
    .B(_0581_),
    .Y(_0137_));
 sg13g2_nand2_2 _2412_ (.Y(_0582_),
    .A(\simon1.state[7] ),
    .B(_0794_));
 sg13g2_nor2b_1 _2413_ (.A(net57),
    .B_N(net56),
    .Y(_0583_));
 sg13g2_o21ai_1 _2414_ (.B1(net60),
    .Y(_0584_),
    .A1(_1033_),
    .A2(net43));
 sg13g2_and2_1 _2415_ (.A(_0583_),
    .B(_0584_),
    .X(_0585_));
 sg13g2_nor3_1 _2416_ (.A(_0032_),
    .B(_0582_),
    .C(_0585_),
    .Y(_0586_));
 sg13g2_o21ai_1 _2417_ (.B1(_0853_),
    .Y(_0587_),
    .A1(_0582_),
    .A2(_0585_));
 sg13g2_o21ai_1 _2418_ (.B1(_0587_),
    .Y(_0588_),
    .A1(net43),
    .A2(_0586_));
 sg13g2_nand2b_1 _2419_ (.Y(_0589_),
    .B(_0588_),
    .A_N(_1045_));
 sg13g2_nand3_1 _2420_ (.B(_0853_),
    .C(_1057_),
    .A(_0835_),
    .Y(_0590_));
 sg13g2_nor2_1 _2421_ (.A(\simon1.state[2] ),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_or2_1 _2422_ (.X(_0592_),
    .B(_0591_),
    .A(_0589_));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]));
 sg13g2_nand2b_1 _2425_ (.Y(_0595_),
    .B(net58),
    .A_N(net55));
 sg13g2_nand2_1 _2426_ (.Y(_0596_),
    .A(_1035_),
    .B(_0595_));
 sg13g2_nor2_1 _2427_ (.A(_1069_),
    .B(_0595_),
    .Y(_0597_));
 sg13g2_a21o_1 _2428_ (.A2(_0596_),
    .A1(_1059_),
    .B1(_0597_),
    .X(_0598_));
 sg13g2_a22oi_1 _2429_ (.Y(_0599_),
    .B1(_0598_),
    .B2(net63),
    .A2(_0849_),
    .A1(net59));
 sg13g2_nor3_2 _2430_ (.A(_0582_),
    .B(_1047_),
    .C(_1051_),
    .Y(_0600_));
 sg13g2_nand2b_1 _2431_ (.Y(_0601_),
    .B(_0600_),
    .A_N(\simon1.millis_counter[0] ));
 sg13g2_a21oi_1 _2432_ (.A1(_0599_),
    .A2(_0601_),
    .Y(_0602_),
    .B1(_0589_));
 sg13g2_a21oi_1 _2433_ (.A1(\simon1.play1.freq[0] ),
    .A2(net21),
    .Y(_0603_),
    .B1(_0602_));
 sg13g2_nor2_1 _2434_ (.A(net89),
    .B(_0603_),
    .Y(_0141_));
 sg13g2_nand2b_1 _2435_ (.Y(_0604_),
    .B(_0595_),
    .A_N(_1038_));
 sg13g2_nor2_1 _2436_ (.A(\simon1.user_input[0] ),
    .B(_1026_),
    .Y(_0605_));
 sg13g2_nor2_1 _2437_ (.A(_1022_),
    .B(\simon1.user_input[1] ),
    .Y(_0606_));
 sg13g2_or2_1 _2438_ (.X(_0607_),
    .B(_0606_),
    .A(_0605_));
 sg13g2_nor4_1 _2439_ (.A(\simon1.state[7] ),
    .B(net64),
    .C(net62),
    .D(\simon1.state[6] ),
    .Y(_0608_));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]));
 sg13g2_a221oi_1 _2441_ (.B2(_0869_),
    .C1(net53),
    .B1(_0607_),
    .A1(net64),
    .Y(_0610_),
    .A2(_0604_));
 sg13g2_xor2_1 _2442_ (.B(\simon1.millis_counter[0] ),
    .A(\simon1.millis_counter[1] ),
    .X(_0611_));
 sg13g2_o21ai_1 _2443_ (.B1(_1039_),
    .Y(_0612_),
    .A1(_1051_),
    .A2(_0611_));
 sg13g2_nand2_1 _2444_ (.Y(_0613_),
    .A(_0849_),
    .B(_0612_));
 sg13g2_xnor2_1 _2445_ (.Y(_0614_),
    .A(net44),
    .B(_0830_));
 sg13g2_a221oi_1 _2446_ (.B2(net53),
    .C1(net21),
    .B1(_0614_),
    .A1(_0610_),
    .Y(_0615_),
    .A2(_0613_));
 sg13g2_a21oi_1 _2447_ (.A1(\simon1.play1.freq[1] ),
    .A2(net21),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_nor2_1 _2448_ (.A(net91),
    .B(_0616_),
    .Y(_0142_));
 sg13g2_nor2_1 _2449_ (.A(\simon1.millis_counter[1] ),
    .B(\simon1.millis_counter[0] ),
    .Y(_0617_));
 sg13g2_nor2b_1 _2450_ (.A(_0617_),
    .B_N(\simon1.millis_counter[2] ),
    .Y(_0618_));
 sg13g2_o21ai_1 _2451_ (.B1(net56),
    .Y(_0619_),
    .A1(_1050_),
    .A2(_0618_));
 sg13g2_nand3_1 _2452_ (.B(_1038_),
    .C(_0619_),
    .A(_0849_),
    .Y(_0620_));
 sg13g2_a21oi_1 _2453_ (.A1(_1026_),
    .A2(net41),
    .Y(_0621_),
    .B1(net53));
 sg13g2_nand2_1 _2454_ (.Y(_0622_),
    .A(_0830_),
    .B(net53));
 sg13g2_inv_1 _2455_ (.Y(_0623_),
    .A(_0622_));
 sg13g2_a21oi_1 _2456_ (.A1(_0620_),
    .A2(_0621_),
    .Y(_0624_),
    .B1(_0623_));
 sg13g2_mux2_1 _2457_ (.A0(_0624_),
    .A1(\simon1.play1.freq[2] ),
    .S(net21),
    .X(_0625_));
 sg13g2_and2_1 _2458_ (.A(net96),
    .B(_0625_),
    .X(_0143_));
 sg13g2_nor2b_1 _2459_ (.A(\simon1.play1.freq[3] ),
    .B_N(net21),
    .Y(_0626_));
 sg13g2_xnor2_1 _2460_ (.Y(_0627_),
    .A(_0019_),
    .B(_0618_));
 sg13g2_o21ai_1 _2461_ (.B1(_1039_),
    .Y(_0628_),
    .A1(_1051_),
    .A2(_0627_));
 sg13g2_o21ai_1 _2462_ (.B1(net64),
    .Y(_0629_),
    .A1(net59),
    .A2(_1034_));
 sg13g2_a21oi_1 _2463_ (.A1(net60),
    .A2(net55),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_a221oi_1 _2464_ (.B2(_0849_),
    .C1(_0630_),
    .B1(_0628_),
    .A1(net41),
    .Y(_0631_),
    .A2(_0605_));
 sg13g2_o21ai_1 _2465_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net44),
    .A2(_0622_));
 sg13g2_nor2_1 _2466_ (.A(net21),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_nor3_1 _2467_ (.A(net91),
    .B(_0626_),
    .C(_0633_),
    .Y(_0144_));
 sg13g2_nor2_1 _2468_ (.A(_1022_),
    .B(_1026_),
    .Y(_0634_));
 sg13g2_a221oi_1 _2469_ (.B2(net41),
    .C1(net22),
    .B1(_0634_),
    .A1(net44),
    .Y(_0635_),
    .A2(_0623_));
 sg13g2_nand2_1 _2470_ (.Y(_0636_),
    .A(net60),
    .B(_0583_));
 sg13g2_o21ai_1 _2471_ (.B1(_0636_),
    .Y(_0637_),
    .A1(net60),
    .A2(_0595_));
 sg13g2_nand2b_1 _2472_ (.Y(_0638_),
    .B(_0873_),
    .A_N(_0617_));
 sg13g2_nand2_1 _2473_ (.Y(_0639_),
    .A(_0019_),
    .B(_0638_));
 sg13g2_xor2_1 _2474_ (.B(_0639_),
    .A(_0020_),
    .X(_0640_));
 sg13g2_a22oi_1 _2475_ (.Y(_0641_),
    .B1(_0640_),
    .B2(_0600_),
    .A2(_0637_),
    .A1(net64));
 sg13g2_a221oi_1 _2476_ (.B2(_0641_),
    .C1(net91),
    .B1(_0635_),
    .A1(_0235_),
    .Y(_0145_),
    .A2(net22));
 sg13g2_nor3_1 _2477_ (.A(\simon1.millis_counter[4] ),
    .B(\simon1.millis_counter[3] ),
    .C(_0618_),
    .Y(_0642_));
 sg13g2_nor2_1 _2478_ (.A(_1047_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nand4_1 _2479_ (.B(_1060_),
    .C(_0794_),
    .A(_1059_),
    .Y(_0644_),
    .D(_0590_));
 sg13g2_nor3_1 _2480_ (.A(net21),
    .B(_0643_),
    .C(_0644_),
    .Y(_0645_));
 sg13g2_a21oi_1 _2481_ (.A1(net81),
    .A2(net22),
    .Y(_0646_),
    .B1(_0645_));
 sg13g2_nor2_1 _2482_ (.A(net91),
    .B(_0646_),
    .Y(_0146_));
 sg13g2_a21o_1 _2483_ (.A2(_0032_),
    .A1(net56),
    .B1(_1038_),
    .X(_0647_));
 sg13g2_a21oi_1 _2484_ (.A1(net64),
    .A2(_0647_),
    .Y(_0648_),
    .B1(net53));
 sg13g2_nor2_1 _2485_ (.A(_0582_),
    .B(_0643_),
    .Y(_0649_));
 sg13g2_a22oi_1 _2486_ (.Y(_0650_),
    .B1(_0649_),
    .B2(_1034_),
    .A2(net41),
    .A1(_1022_));
 sg13g2_a22oi_1 _2487_ (.Y(_0651_),
    .B1(_0648_),
    .B2(_0650_),
    .A2(net53),
    .A1(net44));
 sg13g2_mux2_1 _2488_ (.A0(_0651_),
    .A1(net80),
    .S(net22),
    .X(_0652_));
 sg13g2_and2_1 _2489_ (.A(net97),
    .B(_0652_),
    .X(_0147_));
 sg13g2_xnor2_1 _2490_ (.Y(_0653_),
    .A(net59),
    .B(net57));
 sg13g2_nor3_1 _2491_ (.A(net55),
    .B(_0912_),
    .C(_0653_),
    .Y(_0654_));
 sg13g2_nor2_1 _2492_ (.A(_0608_),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_nor2_1 _2493_ (.A(_0582_),
    .B(_1047_),
    .Y(_0656_));
 sg13g2_nor2_1 _2494_ (.A(\simon1.user_input[0] ),
    .B(\simon1.user_input[1] ),
    .Y(_0657_));
 sg13g2_a22oi_1 _2495_ (.Y(_0658_),
    .B1(_0657_),
    .B2(net41),
    .A2(_0642_),
    .A1(_0656_));
 sg13g2_a221oi_1 _2496_ (.B2(_0658_),
    .C1(_0623_),
    .B1(_0655_),
    .A1(net44),
    .Y(_0659_),
    .A2(net53));
 sg13g2_mux2_1 _2497_ (.A0(_0659_),
    .A1(\simon1.play1.freq[7] ),
    .S(net22),
    .X(_0660_));
 sg13g2_and2_1 _2498_ (.A(net1),
    .B(_0660_),
    .X(_0148_));
 sg13g2_and2_1 _2499_ (.A(_0329_),
    .B(net22),
    .X(_0661_));
 sg13g2_nand2_1 _2500_ (.Y(_0662_),
    .A(_0816_),
    .B(net53));
 sg13g2_o21ai_1 _2501_ (.B1(net55),
    .Y(_0663_),
    .A1(_1059_),
    .A2(_0032_));
 sg13g2_a221oi_1 _2502_ (.B2(net57),
    .C1(_0912_),
    .B1(_0663_),
    .A1(net55),
    .Y(_0664_),
    .A2(_0034_));
 sg13g2_nor2b_1 _2503_ (.A(_0657_),
    .B_N(net41),
    .Y(_0665_));
 sg13g2_nor2_1 _2504_ (.A(_0664_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_nand4_1 _2505_ (.B(_0020_),
    .C(_0600_),
    .A(_0019_),
    .Y(_0667_),
    .D(_0638_));
 sg13g2_nand4_1 _2506_ (.B(_0662_),
    .C(_0666_),
    .A(_0622_),
    .Y(_0668_),
    .D(_0667_));
 sg13g2_nor2_1 _2507_ (.A(net22),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_nor3_1 _2508_ (.A(net92),
    .B(_0661_),
    .C(_0669_),
    .Y(_0149_));
 sg13g2_o21ai_1 _2509_ (.B1(_1039_),
    .Y(_0670_),
    .A1(_1051_),
    .A2(_0642_));
 sg13g2_a22oi_1 _2510_ (.Y(_0671_),
    .B1(_0670_),
    .B2(_0849_),
    .A2(_0596_),
    .A1(net64));
 sg13g2_a221oi_1 _2511_ (.B2(_0671_),
    .C1(net91),
    .B1(_0635_),
    .A1(_0346_),
    .Y(_0150_),
    .A2(net21));
 sg13g2_o21ai_1 _2512_ (.B1(_0849_),
    .Y(_0672_),
    .A1(net43),
    .A2(_1039_));
 sg13g2_a21oi_1 _2513_ (.A1(\simon1.state[0] ),
    .A2(_0794_),
    .Y(_0673_),
    .B1(_0859_));
 sg13g2_nor4_1 _2514_ (.A(\simon1.state[0] ),
    .B(\simon1.state[2] ),
    .C(\simon1.state[1] ),
    .D(_0590_),
    .Y(_0674_));
 sg13g2_nor3_1 _2515_ (.A(net41),
    .B(_1045_),
    .C(_0674_),
    .Y(_0675_));
 sg13g2_nand3_1 _2516_ (.B(_0673_),
    .C(_0675_),
    .A(_0672_),
    .Y(_0676_));
 sg13g2_o21ai_1 _2517_ (.B1(_0853_),
    .Y(_0677_),
    .A1(_0835_),
    .A2(_0833_));
 sg13g2_nor2b_1 _2518_ (.A(_0908_),
    .B_N(_0677_),
    .Y(_0678_));
 sg13g2_o21ai_1 _2519_ (.B1(net96),
    .Y(_0679_),
    .A1(_0676_),
    .A2(_0678_));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_xnor2_1 _2521_ (.Y(_0681_),
    .A(\simon1.millis_counter[0] ),
    .B(_1159_));
 sg13g2_nor2_1 _2522_ (.A(net23),
    .B(_0681_),
    .Y(_0151_));
 sg13g2_nand2_1 _2523_ (.Y(_0682_),
    .A(_1159_),
    .B(_0611_));
 sg13g2_or2_1 _2524_ (.X(_0683_),
    .B(_1159_),
    .A(_0017_));
 sg13g2_a21oi_1 _2525_ (.A1(_0682_),
    .A2(_0683_),
    .Y(_0152_),
    .B1(net23));
 sg13g2_and3_1 _2526_ (.X(_0684_),
    .A(\simon1.millis_counter[1] ),
    .B(\simon1.millis_counter[0] ),
    .C(_1159_));
 sg13g2_xor2_1 _2527_ (.B(_0684_),
    .A(_0018_),
    .X(_0685_));
 sg13g2_nor2_1 _2528_ (.A(net23),
    .B(_0685_),
    .Y(_0153_));
 sg13g2_nand2_1 _2529_ (.Y(_0686_),
    .A(\simon1.millis_counter[2] ),
    .B(_0684_));
 sg13g2_xnor2_1 _2530_ (.Y(_0687_),
    .A(_0019_),
    .B(_0686_));
 sg13g2_nor2_1 _2531_ (.A(net23),
    .B(_0687_),
    .Y(_0154_));
 sg13g2_and3_1 _2532_ (.X(_0688_),
    .A(\simon1.millis_counter[2] ),
    .B(\simon1.millis_counter[3] ),
    .C(_0684_));
 sg13g2_xor2_1 _2533_ (.B(_0688_),
    .A(_0020_),
    .X(_0689_));
 sg13g2_nor2_1 _2534_ (.A(net23),
    .B(_0689_),
    .Y(_0155_));
 sg13g2_and2_1 _2535_ (.A(\simon1.millis_counter[4] ),
    .B(_0688_),
    .X(_0690_));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[4]));
 sg13g2_xor2_1 _2537_ (.B(_0690_),
    .A(_0021_),
    .X(_0692_));
 sg13g2_nor2_1 _2538_ (.A(_0679_),
    .B(_0692_),
    .Y(_0156_));
 sg13g2_nand2_1 _2539_ (.Y(_0693_),
    .A(\simon1.millis_counter[5] ),
    .B(_0690_));
 sg13g2_xnor2_1 _2540_ (.Y(_0694_),
    .A(_0022_),
    .B(_0693_));
 sg13g2_nor2_1 _2541_ (.A(_0679_),
    .B(_0694_),
    .Y(_0157_));
 sg13g2_nand3_1 _2542_ (.B(\simon1.millis_counter[6] ),
    .C(_0690_),
    .A(\simon1.millis_counter[5] ),
    .Y(_0695_));
 sg13g2_xnor2_1 _2543_ (.Y(_0696_),
    .A(_0023_),
    .B(_0695_));
 sg13g2_nor2_1 _2544_ (.A(net23),
    .B(_0696_),
    .Y(_0158_));
 sg13g2_and2_1 _2545_ (.A(_0875_),
    .B(_0690_),
    .X(_0697_));
 sg13g2_xor2_1 _2546_ (.B(_0697_),
    .A(_0024_),
    .X(_0698_));
 sg13g2_nor2_1 _2547_ (.A(net23),
    .B(_0698_),
    .Y(_0159_));
 sg13g2_nand2_1 _2548_ (.Y(_0699_),
    .A(\simon1.millis_counter[8] ),
    .B(_0697_));
 sg13g2_xnor2_1 _2549_ (.Y(_0700_),
    .A(_0025_),
    .B(_0699_));
 sg13g2_nor2_1 _2550_ (.A(net23),
    .B(_0700_),
    .Y(_0160_));
 sg13g2_nor2_2 _2551_ (.A(net61),
    .B(\simon1.state[4] ),
    .Y(_0701_));
 sg13g2_nor2_1 _2552_ (.A(_0031_),
    .B(_0908_),
    .Y(_0702_));
 sg13g2_mux2_1 _2553_ (.A0(net61),
    .A1(_0702_),
    .S(_1196_),
    .X(_0703_));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_nor2_1 _2555_ (.A(_0701_),
    .B(_0703_),
    .Y(_0705_));
 sg13g2_nand2_1 _2556_ (.Y(_0706_),
    .A(net61),
    .B(net70));
 sg13g2_nand2_1 _2557_ (.Y(_0707_),
    .A(_0705_),
    .B(_0706_));
 sg13g2_o21ai_1 _2558_ (.B1(net70),
    .Y(_0708_),
    .A1(_0701_),
    .A2(_0703_));
 sg13g2_a21oi_1 _2559_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0177_),
    .B1(net86));
 sg13g2_a21oi_1 _2560_ (.A1(net70),
    .A2(_1196_),
    .Y(_0709_),
    .B1(_0835_));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_o21ai_1 _2562_ (.B1(\simon1.seq_length[1] ),
    .Y(_0711_),
    .A1(_0701_),
    .A2(_0709_));
 sg13g2_nor3_1 _2563_ (.A(\simon1.seq_length[1] ),
    .B(_0702_),
    .C(_0706_),
    .Y(_0712_));
 sg13g2_and2_1 _2564_ (.A(\simon1.seq_length[1] ),
    .B(_0702_),
    .X(_0713_));
 sg13g2_o21ai_1 _2565_ (.B1(_1196_),
    .Y(_0714_),
    .A1(_0712_),
    .A2(_0713_));
 sg13g2_a21oi_1 _2566_ (.A1(_0711_),
    .A2(_0714_),
    .Y(_0178_),
    .B1(net86));
 sg13g2_o21ai_1 _2567_ (.B1(\simon1.seq_length[2] ),
    .Y(_0715_),
    .A1(_0701_),
    .A2(_0703_));
 sg13g2_nand2_1 _2568_ (.Y(_0716_),
    .A(net70),
    .B(\simon1.seq_length[1] ));
 sg13g2_xnor2_1 _2569_ (.Y(_0717_),
    .A(_0889_),
    .B(_0716_));
 sg13g2_nand3_1 _2570_ (.B(_0705_),
    .C(_0717_),
    .A(net61),
    .Y(_0718_));
 sg13g2_a21oi_1 _2571_ (.A1(_0715_),
    .A2(_0718_),
    .Y(_0179_),
    .B1(net86));
 sg13g2_o21ai_1 _2572_ (.B1(net66),
    .Y(_0719_),
    .A1(_0701_),
    .A2(_0703_));
 sg13g2_nand3_1 _2573_ (.B(net67),
    .C(\simon1.seq_length[1] ),
    .A(net70),
    .Y(_0720_));
 sg13g2_xor2_1 _2574_ (.B(_0720_),
    .A(_0029_),
    .X(_0721_));
 sg13g2_nand3_1 _2575_ (.B(_0705_),
    .C(_0721_),
    .A(net61),
    .Y(_0722_));
 sg13g2_a21oi_1 _2576_ (.A1(_0719_),
    .A2(_0722_),
    .Y(_0180_),
    .B1(net87));
 sg13g2_o21ai_1 _2577_ (.B1(\simon1.seq_length[4] ),
    .Y(_0723_),
    .A1(_0701_),
    .A2(_0703_));
 sg13g2_nand4_1 _2578_ (.B(net67),
    .C(net66),
    .A(net70),
    .Y(_0724_),
    .D(\simon1.seq_length[1] ));
 sg13g2_xor2_1 _2579_ (.B(_0724_),
    .A(_0030_),
    .X(_0725_));
 sg13g2_nand3_1 _2580_ (.B(_0705_),
    .C(_0725_),
    .A(net61),
    .Y(_0726_));
 sg13g2_a21oi_1 _2581_ (.A1(_0723_),
    .A2(_0726_),
    .Y(_0181_),
    .B1(net87));
 sg13g2_nor4_2 _2582_ (.A(\simon1.state[2] ),
    .B(\simon1.state[1] ),
    .C(_0848_),
    .Y(_0727_),
    .D(_0590_));
 sg13g2_a21oi_2 _2583_ (.B1(\simon1.state[4] ),
    .Y(_0728_),
    .A2(_0843_),
    .A1(\simon1.state[6] ));
 sg13g2_o21ai_1 _2584_ (.B1(_0728_),
    .Y(_0729_),
    .A1(_0855_),
    .A2(_0582_));
 sg13g2_a221oi_1 _2585_ (.B2(_0915_),
    .C1(_0729_),
    .B1(_0727_),
    .A1(net62),
    .Y(_0730_),
    .A2(_0657_));
 sg13g2_nand2_1 _2586_ (.Y(_0731_),
    .A(_0835_),
    .B(\simon1.state[2] ));
 sg13g2_nor2_1 _2587_ (.A(net44),
    .B(_0731_),
    .Y(_0732_));
 sg13g2_nand2b_1 _2588_ (.Y(_0733_),
    .B(_0732_),
    .A_N(_0830_));
 sg13g2_o21ai_1 _2589_ (.B1(net97),
    .Y(_0734_),
    .A1(net14),
    .A2(_0728_));
 sg13g2_a21oi_1 _2590_ (.A1(_0730_),
    .A2(_0733_),
    .Y(_0182_),
    .B1(_0734_));
 sg13g2_nor2b_1 _2591_ (.A(_0731_),
    .B_N(net44),
    .Y(_0735_));
 sg13g2_nand2b_1 _2592_ (.Y(_0736_),
    .B(_0735_),
    .A_N(_0830_));
 sg13g2_a221oi_1 _2593_ (.B2(_0839_),
    .C1(_0729_),
    .B1(_0727_),
    .A1(net62),
    .Y(_0737_),
    .A2(_0606_));
 sg13g2_o21ai_1 _2594_ (.B1(net97),
    .Y(_0738_),
    .A1(net15),
    .A2(_0728_));
 sg13g2_a21oi_1 _2595_ (.A1(_0736_),
    .A2(_0737_),
    .Y(_0183_),
    .B1(_0738_));
 sg13g2_nand2b_1 _2596_ (.Y(_0739_),
    .B(\simon1.millis_counter[9] ),
    .A_N(\simon1.millis_counter[8] ));
 sg13g2_a221oi_1 _2597_ (.B2(_0739_),
    .C1(_0729_),
    .B1(_0727_),
    .A1(net62),
    .Y(_0740_),
    .A2(_0605_));
 sg13g2_nand2_1 _2598_ (.Y(_0741_),
    .A(_0830_),
    .B(_0732_));
 sg13g2_o21ai_1 _2599_ (.B1(net97),
    .Y(_0742_),
    .A1(net16),
    .A2(_0728_));
 sg13g2_a21oi_1 _2600_ (.A1(_0740_),
    .A2(_0741_),
    .Y(_0184_),
    .B1(_0742_));
 sg13g2_a221oi_1 _2601_ (.B2(_1048_),
    .C1(_0729_),
    .B1(_0727_),
    .A1(net62),
    .Y(_0743_),
    .A2(_0634_));
 sg13g2_nand2_1 _2602_ (.Y(_0744_),
    .A(_0830_),
    .B(_0735_));
 sg13g2_o21ai_1 _2603_ (.B1(net97),
    .Y(_0745_),
    .A1(net17),
    .A2(_0728_));
 sg13g2_a21oi_1 _2604_ (.A1(_0743_),
    .A2(_0744_),
    .Y(_0185_),
    .B1(_0745_));
 sg13g2_dfrbp_1 _2605_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net102),
    .D(_0082_),
    .Q_N(_1339_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _2606_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_0083_),
    .Q_N(_1338_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _2607_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net104),
    .D(_0084_),
    .Q_N(_1337_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _2608_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net105),
    .D(_0085_),
    .Q_N(_1336_),
    .Q(_0003_));
 sg13g2_dfrbp_1 _2609_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net106),
    .D(_0086_),
    .Q_N(_1335_),
    .Q(_0004_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi ttsimon_101 (.L_HI(net101));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 _2613_ (.A(net107),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2614_ (.A(net108),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2615_ (.A(net109),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2616_ (.A(net110),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2617_ (.A(net111),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2618_ (.A(net112),
    .X(uio_oe[6]));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 _2620_ (.A(net99),
    .X(uio_out[7]));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 _2622_ (.A(net100),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \simon1.millis_counter[0]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net113),
    .D(_0151_),
    .Q_N(_1276_),
    .Q(\simon1.millis_counter[0] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[1]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net114),
    .D(_0152_),
    .Q_N(_0017_),
    .Q(\simon1.millis_counter[1] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[2]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net115),
    .D(_0153_),
    .Q_N(_0018_),
    .Q(\simon1.millis_counter[2] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[3]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net116),
    .D(_0154_),
    .Q_N(_0019_),
    .Q(\simon1.millis_counter[3] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[4]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net117),
    .D(_0155_),
    .Q_N(_0020_),
    .Q(\simon1.millis_counter[4] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[5]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net118),
    .D(_0156_),
    .Q_N(_0021_),
    .Q(\simon1.millis_counter[5] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[6]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net119),
    .D(_0157_),
    .Q_N(_0022_),
    .Q(\simon1.millis_counter[6] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[7]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net120),
    .D(_0158_),
    .Q_N(_0023_),
    .Q(\simon1.millis_counter[7] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[8]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net121),
    .D(_0159_),
    .Q_N(_0024_),
    .Q(\simon1.millis_counter[8] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[9]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net122),
    .D(_0160_),
    .Q_N(_0025_),
    .Q(\simon1.millis_counter[9] ));
 sg13g2_dfrbp_1 \simon1.next_random[0]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net123),
    .D(_0136_),
    .Q_N(_0037_),
    .Q(\simon1.next_random[0] ));
 sg13g2_dfrbp_1 \simon1.next_random[1]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net124),
    .D(_0137_),
    .Q_N(_1288_),
    .Q(\simon1.next_random[1] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[0]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net125),
    .D(_0141_),
    .Q_N(_1286_),
    .Q(\simon1.play1.freq[0] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[1]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net126),
    .D(_0142_),
    .Q_N(_1285_),
    .Q(\simon1.play1.freq[1] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[2]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net127),
    .D(_0143_),
    .Q_N(_1284_),
    .Q(\simon1.play1.freq[2] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[3]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net128),
    .D(_0144_),
    .Q_N(_1283_),
    .Q(\simon1.play1.freq[3] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[4]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net129),
    .D(_0145_),
    .Q_N(_1282_),
    .Q(\simon1.play1.freq[4] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[5]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net130),
    .D(_0146_),
    .Q_N(_1281_),
    .Q(\simon1.play1.freq[5] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[6]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net131),
    .D(_0147_),
    .Q_N(_1280_),
    .Q(\simon1.play1.freq[6] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[7]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net132),
    .D(_0148_),
    .Q_N(_1279_),
    .Q(\simon1.play1.freq[7] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[8]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net133),
    .D(_0149_),
    .Q_N(_1278_),
    .Q(\simon1.play1.freq[8] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[9]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net134),
    .D(_0150_),
    .Q_N(_1277_),
    .Q(\simon1.play1.freq[9] ));
 sg13g2_dfrbp_1 \simon1.play1.sound$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net135),
    .D(_0130_),
    .Q_N(_0013_),
    .Q(net18));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[0]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(_0098_),
    .Q_N(_1323_),
    .Q(\simon1.play1.tick_counter[0] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[10]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net137),
    .D(_0108_),
    .Q_N(_0035_),
    .Q(\simon1.play1.tick_counter[10] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[11]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net138),
    .D(_0109_),
    .Q_N(_1313_),
    .Q(\simon1.play1.tick_counter[11] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[12]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net139),
    .D(_0110_),
    .Q_N(_1312_),
    .Q(\simon1.play1.tick_counter[12] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[13]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net140),
    .D(_0111_),
    .Q_N(_1311_),
    .Q(\simon1.play1.tick_counter[13] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[14]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net141),
    .D(_0112_),
    .Q_N(_1310_),
    .Q(\simon1.play1.tick_counter[14] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[15]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net142),
    .D(_0113_),
    .Q_N(_1309_),
    .Q(\simon1.play1.tick_counter[15] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[16]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net143),
    .D(_0114_),
    .Q_N(_1308_),
    .Q(\simon1.play1.tick_counter[16] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[17]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net144),
    .D(_0115_),
    .Q_N(_1307_),
    .Q(\simon1.play1.tick_counter[17] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[18]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net145),
    .D(_0116_),
    .Q_N(_1306_),
    .Q(\simon1.play1.tick_counter[18] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[19]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net146),
    .D(_0117_),
    .Q_N(_1305_),
    .Q(\simon1.play1.tick_counter[19] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[1]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net147),
    .D(_0099_),
    .Q_N(_1322_),
    .Q(\simon1.play1.tick_counter[1] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[20]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net148),
    .D(_0118_),
    .Q_N(_1304_),
    .Q(\simon1.play1.tick_counter[20] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[21]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net149),
    .D(_0119_),
    .Q_N(_1303_),
    .Q(\simon1.play1.tick_counter[21] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[22]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net150),
    .D(_0120_),
    .Q_N(_1302_),
    .Q(\simon1.play1.tick_counter[22] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[23]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net151),
    .D(_0121_),
    .Q_N(_1301_),
    .Q(\simon1.play1.tick_counter[23] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[24]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net152),
    .D(_0122_),
    .Q_N(_1300_),
    .Q(\simon1.play1.tick_counter[24] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[25]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net153),
    .D(_0123_),
    .Q_N(_1299_),
    .Q(\simon1.play1.tick_counter[25] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[26]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net154),
    .D(_0124_),
    .Q_N(_1298_),
    .Q(\simon1.play1.tick_counter[26] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[27]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net155),
    .D(_0125_),
    .Q_N(_1297_),
    .Q(\simon1.play1.tick_counter[27] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[28]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net156),
    .D(_0126_),
    .Q_N(_1296_),
    .Q(\simon1.play1.tick_counter[28] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[29]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net157),
    .D(_0127_),
    .Q_N(_1295_),
    .Q(\simon1.play1.tick_counter[29] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[2]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net158),
    .D(_0100_),
    .Q_N(_1321_),
    .Q(\simon1.play1.tick_counter[2] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[30]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net159),
    .D(_0128_),
    .Q_N(_1294_),
    .Q(\simon1.play1.tick_counter[30] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[31]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net160),
    .D(_0129_),
    .Q_N(_1293_),
    .Q(\simon1.play1.tick_counter[31] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[3]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net161),
    .D(_0101_),
    .Q_N(_1320_),
    .Q(\simon1.play1.tick_counter[3] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[4]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net162),
    .D(_0102_),
    .Q_N(_1319_),
    .Q(\simon1.play1.tick_counter[4] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[5]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net163),
    .D(_0103_),
    .Q_N(_1318_),
    .Q(\simon1.play1.tick_counter[5] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[6]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net164),
    .D(_0104_),
    .Q_N(_1317_),
    .Q(\simon1.play1.tick_counter[6] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[7]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net165),
    .D(_0105_),
    .Q_N(_1316_),
    .Q(\simon1.play1.tick_counter[7] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[8]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net166),
    .D(_0106_),
    .Q_N(_1315_),
    .Q(\simon1.play1.tick_counter[8] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[9]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net167),
    .D(_0107_),
    .Q_N(_1314_),
    .Q(\simon1.play1.tick_counter[9] ));
 sg13g2_dfrbp_1 \simon1.score1.active_digit$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net168),
    .D(_0081_),
    .Q_N(_0016_),
    .Q(\simon1.score1.active_digit ));
 sg13g2_dfrbp_1 \simon1.score1.ena$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net169),
    .D(_0132_),
    .Q_N(_0026_),
    .Q(\simon1.score1.ena ));
 sg13g2_dfrbp_1 \simon1.score1.inc$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net170),
    .D(_0133_),
    .Q_N(_1291_),
    .Q(\simon1.score1.inc ));
 sg13g2_dfrbp_1 \simon1.score1.ones[0]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net171),
    .D(_0090_),
    .Q_N(_1331_),
    .Q(\simon1.score1.ones[0] ));
 sg13g2_dfrbp_1 \simon1.score1.ones[1]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net172),
    .D(_0091_),
    .Q_N(_1330_),
    .Q(\simon1.score1.ones[1] ));
 sg13g2_dfrbp_1 \simon1.score1.ones[2]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net173),
    .D(_0092_),
    .Q_N(_1329_),
    .Q(\simon1.score1.ones[2] ));
 sg13g2_dfrbp_1 \simon1.score1.ones[3]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net174),
    .D(_0093_),
    .Q_N(_1328_),
    .Q(\simon1.score1.ones[3] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[0]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net175),
    .D(_0094_),
    .Q_N(_1327_),
    .Q(\simon1.score1.tens[0] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[1]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net176),
    .D(_0095_),
    .Q_N(_1326_),
    .Q(\simon1.score1.tens[1] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[2]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net177),
    .D(_0096_),
    .Q_N(_1325_),
    .Q(\simon1.score1.tens[2] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[3]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net178),
    .D(_0097_),
    .Q_N(_1324_),
    .Q(\simon1.score1.tens[3] ));
 sg13g2_dfrbp_1 \simon1.score_rst$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net179),
    .D(_0089_),
    .Q_N(_1332_),
    .Q(\simon1.score_rst ));
 sg13g2_dfrbp_1 \simon1.seq[0][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net180),
    .D(_0038_),
    .Q_N(_1381_),
    .Q(\simon1.seq[0][0] ));
 sg13g2_dfrbp_1 \simon1.seq[0][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net181),
    .D(_0203_),
    .Q_N(_1233_),
    .Q(\simon1.seq[0][1] ));
 sg13g2_dfrbp_1 \simon1.seq[10][0]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net182),
    .D(_0197_),
    .Q_N(_1239_),
    .Q(\simon1.seq[10][0] ));
 sg13g2_dfrbp_1 \simon1.seq[10][1]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net183),
    .D(_0064_),
    .Q_N(_1355_),
    .Q(\simon1.seq[10][1] ));
 sg13g2_dfrbp_1 \simon1.seq[11][0]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net184),
    .D(_0066_),
    .Q_N(_1353_),
    .Q(\simon1.seq[11][0] ));
 sg13g2_dfrbp_1 \simon1.seq[11][1]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net185),
    .D(_0054_),
    .Q_N(_1365_),
    .Q(\simon1.seq[11][1] ));
 sg13g2_dfrbp_1 \simon1.seq[12][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net186),
    .D(_0065_),
    .Q_N(_1354_),
    .Q(\simon1.seq[12][0] ));
 sg13g2_dfrbp_1 \simon1.seq[12][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net187),
    .D(_0042_),
    .Q_N(_1377_),
    .Q(\simon1.seq[12][1] ));
 sg13g2_dfrbp_1 \simon1.seq[13][0]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net188),
    .D(_0063_),
    .Q_N(_1356_),
    .Q(\simon1.seq[13][0] ));
 sg13g2_dfrbp_1 \simon1.seq[13][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net189),
    .D(_0041_),
    .Q_N(_1378_),
    .Q(\simon1.seq[13][1] ));
 sg13g2_dfrbp_1 \simon1.seq[14][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net190),
    .D(_0062_),
    .Q_N(_1357_),
    .Q(\simon1.seq[14][0] ));
 sg13g2_dfrbp_1 \simon1.seq[14][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net191),
    .D(_0040_),
    .Q_N(_1379_),
    .Q(\simon1.seq[14][1] ));
 sg13g2_dfrbp_1 \simon1.seq[15][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net192),
    .D(_0061_),
    .Q_N(_1358_),
    .Q(\simon1.seq[15][0] ));
 sg13g2_dfrbp_1 \simon1.seq[15][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net193),
    .D(_0201_),
    .Q_N(_1235_),
    .Q(\simon1.seq[15][1] ));
 sg13g2_dfrbp_1 \simon1.seq[16][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net194),
    .D(_0060_),
    .Q_N(_1359_),
    .Q(\simon1.seq[16][0] ));
 sg13g2_dfrbp_1 \simon1.seq[16][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net195),
    .D(_0198_),
    .Q_N(_1238_),
    .Q(\simon1.seq[16][1] ));
 sg13g2_dfrbp_1 \simon1.seq[17][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net196),
    .D(_0059_),
    .Q_N(_1360_),
    .Q(\simon1.seq[17][0] ));
 sg13g2_dfrbp_1 \simon1.seq[17][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net197),
    .D(_0196_),
    .Q_N(_1240_),
    .Q(\simon1.seq[17][1] ));
 sg13g2_dfrbp_1 \simon1.seq[18][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net198),
    .D(_0058_),
    .Q_N(_1361_),
    .Q(\simon1.seq[18][0] ));
 sg13g2_dfrbp_1 \simon1.seq[18][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net199),
    .D(_0187_),
    .Q_N(_1249_),
    .Q(\simon1.seq[18][1] ));
 sg13g2_dfrbp_1 \simon1.seq[19][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net200),
    .D(_0057_),
    .Q_N(_1362_),
    .Q(\simon1.seq[19][0] ));
 sg13g2_dfrbp_1 \simon1.seq[19][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net201),
    .D(_0195_),
    .Q_N(_1241_),
    .Q(\simon1.seq[19][1] ));
 sg13g2_dfrbp_1 \simon1.seq[1][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net202),
    .D(_0056_),
    .Q_N(_1363_),
    .Q(\simon1.seq[1][0] ));
 sg13g2_dfrbp_1 \simon1.seq[1][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net203),
    .D(_0200_),
    .Q_N(_1236_),
    .Q(\simon1.seq[1][1] ));
 sg13g2_dfrbp_1 \simon1.seq[20][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net204),
    .D(_0199_),
    .Q_N(_1237_),
    .Q(\simon1.seq[20][0] ));
 sg13g2_dfrbp_1 \simon1.seq[20][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net205),
    .D(_0192_),
    .Q_N(_1244_),
    .Q(\simon1.seq[20][1] ));
 sg13g2_dfrbp_1 \simon1.seq[21][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net206),
    .D(_0055_),
    .Q_N(_1364_),
    .Q(\simon1.seq[21][0] ));
 sg13g2_dfrbp_1 \simon1.seq[21][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net207),
    .D(_0193_),
    .Q_N(_1243_),
    .Q(\simon1.seq[21][1] ));
 sg13g2_dfrbp_1 \simon1.seq[22][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net208),
    .D(_0053_),
    .Q_N(_1366_),
    .Q(\simon1.seq[22][0] ));
 sg13g2_dfrbp_1 \simon1.seq[22][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net209),
    .D(_0190_),
    .Q_N(_1246_),
    .Q(\simon1.seq[22][1] ));
 sg13g2_dfrbp_1 \simon1.seq[23][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net210),
    .D(_0052_),
    .Q_N(_1367_),
    .Q(\simon1.seq[23][0] ));
 sg13g2_dfrbp_1 \simon1.seq[23][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net211),
    .D(_0191_),
    .Q_N(_1245_),
    .Q(\simon1.seq[23][1] ));
 sg13g2_dfrbp_1 \simon1.seq[24][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net212),
    .D(_0051_),
    .Q_N(_1368_),
    .Q(\simon1.seq[24][0] ));
 sg13g2_dfrbp_1 \simon1.seq[24][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net213),
    .D(_0194_),
    .Q_N(_1242_),
    .Q(\simon1.seq[24][1] ));
 sg13g2_dfrbp_1 \simon1.seq[25][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net214),
    .D(_0050_),
    .Q_N(_1369_),
    .Q(\simon1.seq[25][0] ));
 sg13g2_dfrbp_1 \simon1.seq[25][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net215),
    .D(_0189_),
    .Q_N(_1247_),
    .Q(\simon1.seq[25][1] ));
 sg13g2_dfrbp_1 \simon1.seq[26][0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net216),
    .D(_0049_),
    .Q_N(_1370_),
    .Q(\simon1.seq[26][0] ));
 sg13g2_dfrbp_1 \simon1.seq[26][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net217),
    .D(_0188_),
    .Q_N(_1248_),
    .Q(\simon1.seq[26][1] ));
 sg13g2_dfrbp_1 \simon1.seq[27][0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net218),
    .D(_0048_),
    .Q_N(_1371_),
    .Q(\simon1.seq[27][0] ));
 sg13g2_dfrbp_1 \simon1.seq[27][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net219),
    .D(_0186_),
    .Q_N(_1250_),
    .Q(\simon1.seq[27][1] ));
 sg13g2_dfrbp_1 \simon1.seq[28][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net220),
    .D(_0047_),
    .Q_N(_1372_),
    .Q(\simon1.seq[28][0] ));
 sg13g2_dfrbp_1 \simon1.seq[28][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net221),
    .D(_0131_),
    .Q_N(_1292_),
    .Q(\simon1.seq[28][1] ));
 sg13g2_dfrbp_1 \simon1.seq[29][0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net222),
    .D(_0046_),
    .Q_N(_1373_),
    .Q(\simon1.seq[29][0] ));
 sg13g2_dfrbp_1 \simon1.seq[29][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net223),
    .D(_0202_),
    .Q_N(_1234_),
    .Q(\simon1.seq[29][1] ));
 sg13g2_dfrbp_1 \simon1.seq[2][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net224),
    .D(_0045_),
    .Q_N(_1374_),
    .Q(\simon1.seq[2][0] ));
 sg13g2_dfrbp_1 \simon1.seq[2][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net225),
    .D(_0088_),
    .Q_N(_1389_),
    .Q(\simon1.seq[2][1] ));
 sg13g2_dfrbp_1 \simon1.seq[30][0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net226),
    .D(_0080_),
    .Q_N(_1340_),
    .Q(\simon1.seq[30][0] ));
 sg13g2_dfrbp_1 \simon1.seq[30][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net227),
    .D(_0087_),
    .Q_N(_1334_),
    .Q(\simon1.seq[30][1] ));
 sg13g2_dfrbp_1 \simon1.seq[31][0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net228),
    .D(_0044_),
    .Q_N(_1375_),
    .Q(\simon1.seq[31][0] ));
 sg13g2_dfrbp_1 \simon1.seq[31][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net229),
    .D(_0077_),
    .Q_N(_1343_),
    .Q(\simon1.seq[31][1] ));
 sg13g2_dfrbp_1 \simon1.seq[3][0]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net230),
    .D(_0043_),
    .Q_N(_1376_),
    .Q(\simon1.seq[3][0] ));
 sg13g2_dfrbp_1 \simon1.seq[3][1]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net231),
    .D(_0078_),
    .Q_N(_1342_),
    .Q(\simon1.seq[3][1] ));
 sg13g2_dfrbp_1 \simon1.seq[4][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net232),
    .D(_0079_),
    .Q_N(_1341_),
    .Q(\simon1.seq[4][0] ));
 sg13g2_dfrbp_1 \simon1.seq[4][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net233),
    .D(_0076_),
    .Q_N(_1344_),
    .Q(\simon1.seq[4][1] ));
 sg13g2_dfrbp_1 \simon1.seq[5][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net234),
    .D(_0075_),
    .Q_N(_1345_),
    .Q(\simon1.seq[5][0] ));
 sg13g2_dfrbp_1 \simon1.seq[5][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net235),
    .D(_0071_),
    .Q_N(_1349_),
    .Q(\simon1.seq[5][1] ));
 sg13g2_dfrbp_1 \simon1.seq[6][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net236),
    .D(_0074_),
    .Q_N(_1346_),
    .Q(\simon1.seq[6][0] ));
 sg13g2_dfrbp_1 \simon1.seq[6][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net237),
    .D(_0070_),
    .Q_N(_1350_),
    .Q(\simon1.seq[6][1] ));
 sg13g2_dfrbp_1 \simon1.seq[7][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net238),
    .D(_0073_),
    .Q_N(_1347_),
    .Q(\simon1.seq[7][0] ));
 sg13g2_dfrbp_1 \simon1.seq[7][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net239),
    .D(_0069_),
    .Q_N(_1351_),
    .Q(\simon1.seq[7][1] ));
 sg13g2_dfrbp_1 \simon1.seq[8][0]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net240),
    .D(_0072_),
    .Q_N(_1348_),
    .Q(\simon1.seq[8][0] ));
 sg13g2_dfrbp_1 \simon1.seq[8][1]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net241),
    .D(_0039_),
    .Q_N(_1380_),
    .Q(\simon1.seq[8][1] ));
 sg13g2_dfrbp_1 \simon1.seq[9][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net242),
    .D(_0068_),
    .Q_N(_1382_),
    .Q(\simon1.seq[9][0] ));
 sg13g2_dfrbp_1 \simon1.seq[9][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net243),
    .D(_0067_),
    .Q_N(_1352_),
    .Q(\simon1.seq[9][1] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net244),
    .D(_0082_),
    .Q_N(_1259_),
    .Q(\simon1.seq_counter[0] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net245),
    .D(_0083_),
    .Q_N(_1258_),
    .Q(\simon1.seq_counter[1] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net246),
    .D(_0084_),
    .Q_N(_1257_),
    .Q(\simon1.seq_counter[2] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net247),
    .D(_0085_),
    .Q_N(_1256_),
    .Q(\simon1.seq_counter[3] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net248),
    .D(_0086_),
    .Q_N(_1255_),
    .Q(\simon1.seq_counter[4] ));
 sg13g2_dfrbp_1 \simon1.seq_length[0]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net249),
    .D(_0177_),
    .Q_N(_1260_),
    .Q(\simon1.seq_length[0] ));
 sg13g2_dfrbp_1 \simon1.seq_length[1]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net250),
    .D(_0178_),
    .Q_N(_0027_),
    .Q(\simon1.seq_length[1] ));
 sg13g2_dfrbp_1 \simon1.seq_length[2]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net251),
    .D(_0179_),
    .Q_N(_0028_),
    .Q(\simon1.seq_length[2] ));
 sg13g2_dfrbp_1 \simon1.seq_length[3]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net252),
    .D(_0180_),
    .Q_N(_0029_),
    .Q(\simon1.seq_length[3] ));
 sg13g2_dfrbp_1 \simon1.seq_length[4]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net253),
    .D(_0181_),
    .Q_N(_0030_),
    .Q(\simon1.seq_length[4] ));
 sg13g2_dfrbp_1 \simon1.state[0]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net254),
    .D(_0005_),
    .Q_N(_1383_),
    .Q(\simon1.state[0] ));
 sg13g2_dfrbp_1 \simon1.state[1]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net255),
    .D(_0006_),
    .Q_N(_1384_),
    .Q(\simon1.state[1] ));
 sg13g2_dfrbp_1 \simon1.state[2]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net256),
    .D(_0007_),
    .Q_N(_1385_),
    .Q(\simon1.state[2] ));
 sg13g2_dfrbp_1 \simon1.state[3]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net257),
    .D(_0008_),
    .Q_N(_1386_),
    .Q(\simon1.state[3] ));
 sg13g2_dfrbp_1 \simon1.state[4]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net258),
    .D(_0009_),
    .Q_N(_1387_),
    .Q(\simon1.state[4] ));
 sg13g2_dfrbp_1 \simon1.state[5]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net259),
    .D(_0010_),
    .Q_N(_0031_),
    .Q(\simon1.state[5] ));
 sg13g2_dfrbp_1 \simon1.state[6]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net260),
    .D(_0011_),
    .Q_N(_1388_),
    .Q(\simon1.state[6] ));
 sg13g2_dfrbp_1 \simon1.state[7]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net261),
    .D(_0012_),
    .Q_N(_0033_),
    .Q(\simon1.state[7] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[0]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net262),
    .D(_0161_),
    .Q_N(_0036_),
    .Q(\simon1.tick_counter[0] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[10]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net263),
    .D(_0171_),
    .Q_N(_1266_),
    .Q(\simon1.tick_counter[10] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[11]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net264),
    .D(_0172_),
    .Q_N(_1265_),
    .Q(\simon1.tick_counter[11] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[12]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net265),
    .D(_0173_),
    .Q_N(_1264_),
    .Q(\simon1.tick_counter[12] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[13]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net266),
    .D(_0174_),
    .Q_N(_1263_),
    .Q(\simon1.tick_counter[13] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[14]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net267),
    .D(_0175_),
    .Q_N(_1262_),
    .Q(\simon1.tick_counter[14] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[15]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net268),
    .D(_0176_),
    .Q_N(_1261_),
    .Q(\simon1.tick_counter[15] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[1]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net269),
    .D(_0162_),
    .Q_N(_1275_),
    .Q(\simon1.tick_counter[1] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[2]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net270),
    .D(_0163_),
    .Q_N(_1274_),
    .Q(\simon1.tick_counter[2] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[3]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net271),
    .D(_0164_),
    .Q_N(_1273_),
    .Q(\simon1.tick_counter[3] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[4]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net272),
    .D(_0165_),
    .Q_N(_1272_),
    .Q(\simon1.tick_counter[4] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[5]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net273),
    .D(_0166_),
    .Q_N(_1271_),
    .Q(\simon1.tick_counter[5] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[6]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net274),
    .D(_0167_),
    .Q_N(_1270_),
    .Q(\simon1.tick_counter[6] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[7]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net275),
    .D(_0168_),
    .Q_N(_1269_),
    .Q(\simon1.tick_counter[7] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[8]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net276),
    .D(_0169_),
    .Q_N(_1268_),
    .Q(\simon1.tick_counter[8] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[9]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net277),
    .D(_0170_),
    .Q_N(_1267_),
    .Q(\simon1.tick_counter[9] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[0]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net278),
    .D(_0138_),
    .Q_N(_0034_),
    .Q(\simon1.tone_sequence_counter[0] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[1]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net279),
    .D(_0139_),
    .Q_N(_1287_),
    .Q(\simon1.tone_sequence_counter[1] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[2]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net280),
    .D(_0140_),
    .Q_N(_0032_),
    .Q(\simon1.tone_sequence_counter[2] ));
 sg13g2_dfrbp_1 \simon1.user_input[0]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net281),
    .D(_0134_),
    .Q_N(_1290_),
    .Q(\simon1.user_input[0] ));
 sg13g2_dfrbp_1 \simon1.user_input[1]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net282),
    .D(_0135_),
    .Q_N(_1289_),
    .Q(\simon1.user_input[1] ));
 sg13g2_dfrbp_1 \uio_out[0]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net283),
    .D(_0204_),
    .Q_N(_1390_),
    .Q(net7));
 sg13g2_dfrbp_1 \uio_out[1]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net284),
    .D(_0205_),
    .Q_N(_1391_),
    .Q(net8));
 sg13g2_dfrbp_1 \uio_out[2]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net285),
    .D(_0206_),
    .Q_N(_1392_),
    .Q(net9));
 sg13g2_dfrbp_1 \uio_out[3]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net286),
    .D(_0207_),
    .Q_N(_1393_),
    .Q(net10));
 sg13g2_dfrbp_1 \uio_out[4]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net287),
    .D(_0208_),
    .Q_N(_1394_),
    .Q(net11));
 sg13g2_dfrbp_1 \uio_out[5]$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net288),
    .D(_0209_),
    .Q_N(_1395_),
    .Q(net12));
 sg13g2_dfrbp_1 \uio_out[6]$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net289),
    .D(_0210_),
    .Q_N(_1396_),
    .Q(net13));
 sg13g2_dfrbp_1 \uo_out[0]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net290),
    .D(_0182_),
    .Q_N(_1254_),
    .Q(net14));
 sg13g2_dfrbp_1 \uo_out[1]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net291),
    .D(_0183_),
    .Q_N(_1253_),
    .Q(net15));
 sg13g2_dfrbp_1 \uo_out[2]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net292),
    .D(_0184_),
    .Q_N(_1252_),
    .Q(net16));
 sg13g2_dfrbp_1 \uo_out[3]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net293),
    .D(_0185_),
    .Q_N(_1251_),
    .Q(net17));
 sg13g2_dfrbp_1 \uo_out[5]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net294),
    .D(_0014_),
    .Q_N(_1397_),
    .Q(net19));
 sg13g2_dfrbp_1 \uo_out[6]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net295),
    .D(_0015_),
    .Q_N(_1333_),
    .Q(net20));
 sg13g2_tiehi \simon1.play1.tick_counter[11]$_SDFFE_PN0N__138  (.L_HI(net138));
 sg13g2_tiehi \simon1.play1.tick_counter[12]$_SDFFE_PN0N__139  (.L_HI(net139));
 sg13g2_tiehi \simon1.play1.tick_counter[13]$_SDFFE_PN0N__140  (.L_HI(net140));
 sg13g2_tiehi \simon1.play1.tick_counter[14]$_SDFFE_PN0N__141  (.L_HI(net141));
 sg13g2_tiehi \simon1.play1.tick_counter[15]$_SDFFE_PN0N__142  (.L_HI(net142));
 sg13g2_tiehi \simon1.play1.tick_counter[16]$_SDFFE_PN0N__143  (.L_HI(net143));
 sg13g2_tiehi \simon1.play1.tick_counter[17]$_SDFFE_PN0N__144  (.L_HI(net144));
 sg13g2_tiehi \simon1.play1.tick_counter[18]$_SDFFE_PN0N__145  (.L_HI(net145));
 sg13g2_tiehi \simon1.play1.tick_counter[19]$_SDFFE_PN0N__146  (.L_HI(net146));
 sg13g2_tiehi \simon1.play1.tick_counter[1]$_SDFFE_PN0N__147  (.L_HI(net147));
 sg13g2_tiehi \simon1.play1.tick_counter[20]$_SDFFE_PN0N__148  (.L_HI(net148));
 sg13g2_tiehi \simon1.play1.tick_counter[21]$_SDFFE_PN0N__149  (.L_HI(net149));
 sg13g2_tiehi \simon1.play1.tick_counter[22]$_SDFFE_PN0N__150  (.L_HI(net150));
 sg13g2_tiehi \simon1.play1.tick_counter[23]$_SDFFE_PN0N__151  (.L_HI(net151));
 sg13g2_tiehi \simon1.play1.tick_counter[24]$_SDFFE_PN0N__152  (.L_HI(net152));
 sg13g2_tiehi \simon1.play1.tick_counter[25]$_SDFFE_PN0N__153  (.L_HI(net153));
 sg13g2_tiehi \simon1.play1.tick_counter[26]$_SDFFE_PN0N__154  (.L_HI(net154));
 sg13g2_tiehi \simon1.play1.tick_counter[27]$_SDFFE_PN0N__155  (.L_HI(net155));
 sg13g2_tiehi \simon1.play1.tick_counter[28]$_SDFFE_PN0N__156  (.L_HI(net156));
 sg13g2_tiehi \simon1.play1.tick_counter[29]$_SDFFE_PN0N__157  (.L_HI(net157));
 sg13g2_tiehi \simon1.play1.tick_counter[2]$_SDFFE_PN0N__158  (.L_HI(net158));
 sg13g2_tiehi \simon1.play1.tick_counter[30]$_SDFFE_PN0N__159  (.L_HI(net159));
 sg13g2_tiehi \simon1.play1.tick_counter[31]$_SDFFE_PN0N__160  (.L_HI(net160));
 sg13g2_tiehi \simon1.play1.tick_counter[3]$_SDFFE_PN0N__161  (.L_HI(net161));
 sg13g2_tiehi \simon1.play1.tick_counter[4]$_SDFFE_PN0N__162  (.L_HI(net162));
 sg13g2_tiehi \simon1.play1.tick_counter[5]$_SDFFE_PN0N__163  (.L_HI(net163));
 sg13g2_tiehi \simon1.play1.tick_counter[6]$_SDFFE_PN0N__164  (.L_HI(net164));
 sg13g2_tiehi \simon1.play1.tick_counter[7]$_SDFFE_PN0N__165  (.L_HI(net165));
 sg13g2_tiehi \simon1.play1.tick_counter[8]$_SDFFE_PN0N__166  (.L_HI(net166));
 sg13g2_tiehi \simon1.play1.tick_counter[9]$_SDFFE_PN0N__167  (.L_HI(net167));
 sg13g2_tiehi \simon1.score1.active_digit$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \simon1.score1.ena$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \simon1.score1.inc$_SDFF_PN0__170  (.L_HI(net170));
 sg13g2_tiehi \simon1.score1.ones[0]$_SDFFE_PP0P__171  (.L_HI(net171));
 sg13g2_tiehi \simon1.score1.ones[1]$_SDFFE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \simon1.score1.ones[2]$_SDFFE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \simon1.score1.ones[3]$_SDFFE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \simon1.score1.tens[0]$_SDFFE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \simon1.score1.tens[1]$_SDFFE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \simon1.score1.tens[2]$_SDFFE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \simon1.score1.tens[3]$_SDFFE_PP0P__178  (.L_HI(net178));
 sg13g2_tiehi \simon1.score_rst$_SDFF_PN0__179  (.L_HI(net179));
 sg13g2_tiehi \simon1.seq[0][0]$_DFFE_PP__180  (.L_HI(net180));
 sg13g2_tiehi \simon1.seq[0][1]$_DFFE_PP__181  (.L_HI(net181));
 sg13g2_tiehi \simon1.seq[10][0]$_DFFE_PP__182  (.L_HI(net182));
 sg13g2_tiehi \simon1.seq[10][1]$_DFFE_PP__183  (.L_HI(net183));
 sg13g2_tiehi \simon1.seq[11][0]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \simon1.seq[11][1]$_DFFE_PP__185  (.L_HI(net185));
 sg13g2_tiehi \simon1.seq[12][0]$_DFFE_PP__186  (.L_HI(net186));
 sg13g2_tiehi \simon1.seq[12][1]$_DFFE_PP__187  (.L_HI(net187));
 sg13g2_tiehi \simon1.seq[13][0]$_DFFE_PP__188  (.L_HI(net188));
 sg13g2_tiehi \simon1.seq[13][1]$_DFFE_PP__189  (.L_HI(net189));
 sg13g2_tiehi \simon1.seq[14][0]$_DFFE_PP__190  (.L_HI(net190));
 sg13g2_tiehi \simon1.seq[14][1]$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \simon1.seq[15][0]$_DFFE_PP__192  (.L_HI(net192));
 sg13g2_tiehi \simon1.seq[15][1]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \simon1.seq[16][0]$_DFFE_PP__194  (.L_HI(net194));
 sg13g2_tiehi \simon1.seq[16][1]$_DFFE_PP__195  (.L_HI(net195));
 sg13g2_tiehi \simon1.seq[17][0]$_DFFE_PP__196  (.L_HI(net196));
 sg13g2_tiehi \simon1.seq[17][1]$_DFFE_PP__197  (.L_HI(net197));
 sg13g2_tiehi \simon1.seq[18][0]$_DFFE_PP__198  (.L_HI(net198));
 sg13g2_tiehi \simon1.seq[18][1]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \simon1.seq[19][0]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \simon1.seq[19][1]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \simon1.seq[1][0]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \simon1.seq[1][1]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \simon1.seq[20][0]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \simon1.seq[20][1]$_DFFE_PP__205  (.L_HI(net205));
 sg13g2_tiehi \simon1.seq[21][0]$_DFFE_PP__206  (.L_HI(net206));
 sg13g2_tiehi \simon1.seq[21][1]$_DFFE_PP__207  (.L_HI(net207));
 sg13g2_tiehi \simon1.seq[22][0]$_DFFE_PP__208  (.L_HI(net208));
 sg13g2_tiehi \simon1.seq[22][1]$_DFFE_PP__209  (.L_HI(net209));
 sg13g2_tiehi \simon1.seq[23][0]$_DFFE_PP__210  (.L_HI(net210));
 sg13g2_tiehi \simon1.seq[23][1]$_DFFE_PP__211  (.L_HI(net211));
 sg13g2_tiehi \simon1.seq[24][0]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \simon1.seq[24][1]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \simon1.seq[25][0]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \simon1.seq[25][1]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \simon1.seq[26][0]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \simon1.seq[26][1]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \simon1.seq[27][0]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \simon1.seq[27][1]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \simon1.seq[28][0]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \simon1.seq[28][1]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \simon1.seq[29][0]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \simon1.seq[29][1]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \simon1.seq[2][0]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \simon1.seq[2][1]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \simon1.seq[30][0]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \simon1.seq[30][1]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \simon1.seq[31][0]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \simon1.seq[31][1]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \simon1.seq[3][0]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \simon1.seq[3][1]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \simon1.seq[4][0]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \simon1.seq[4][1]$_DFFE_PP__233  (.L_HI(net233));
 sg13g2_tiehi \simon1.seq[5][0]$_DFFE_PP__234  (.L_HI(net234));
 sg13g2_tiehi \simon1.seq[5][1]$_DFFE_PP__235  (.L_HI(net235));
 sg13g2_tiehi \simon1.seq[6][0]$_DFFE_PP__236  (.L_HI(net236));
 sg13g2_tiehi \simon1.seq[6][1]$_DFFE_PP__237  (.L_HI(net237));
 sg13g2_tiehi \simon1.seq[7][0]$_DFFE_PP__238  (.L_HI(net238));
 sg13g2_tiehi \simon1.seq[7][1]$_DFFE_PP__239  (.L_HI(net239));
 sg13g2_tiehi \simon1.seq[8][0]$_DFFE_PP__240  (.L_HI(net240));
 sg13g2_tiehi \simon1.seq[8][1]$_DFFE_PP__241  (.L_HI(net241));
 sg13g2_tiehi \simon1.seq[9][0]$_DFFE_PP__242  (.L_HI(net242));
 sg13g2_tiehi \simon1.seq[9][1]$_DFFE_PP__243  (.L_HI(net243));
 sg13g2_tiehi \simon1.seq_counter[0]$_SDFFE_PN0P__244  (.L_HI(net244));
 sg13g2_tiehi \simon1.seq_counter[1]$_SDFFE_PN0P__245  (.L_HI(net245));
 sg13g2_tiehi \simon1.seq_counter[2]$_SDFFE_PN0P__246  (.L_HI(net246));
 sg13g2_tiehi \simon1.seq_counter[3]$_SDFFE_PN0P__247  (.L_HI(net247));
 sg13g2_tiehi \simon1.seq_counter[4]$_SDFFE_PN0P__248  (.L_HI(net248));
 sg13g2_tiehi \simon1.seq_length[0]$_SDFFE_PN0P__249  (.L_HI(net249));
 sg13g2_tiehi \simon1.seq_length[1]$_SDFFE_PN0P__250  (.L_HI(net250));
 sg13g2_tiehi \simon1.seq_length[2]$_SDFFE_PN0P__251  (.L_HI(net251));
 sg13g2_tiehi \simon1.seq_length[3]$_SDFFE_PN0P__252  (.L_HI(net252));
 sg13g2_tiehi \simon1.seq_length[4]$_SDFFE_PN0P__253  (.L_HI(net253));
 sg13g2_tiehi \simon1.state[0]$_DFF_P__254  (.L_HI(net254));
 sg13g2_tiehi \simon1.state[1]$_DFF_P__255  (.L_HI(net255));
 sg13g2_tiehi \simon1.state[2]$_DFF_P__256  (.L_HI(net256));
 sg13g2_tiehi \simon1.state[3]$_DFF_P__257  (.L_HI(net257));
 sg13g2_tiehi \simon1.state[4]$_DFF_P__258  (.L_HI(net258));
 sg13g2_tiehi \simon1.state[5]$_DFF_P__259  (.L_HI(net259));
 sg13g2_tiehi \simon1.state[6]$_DFF_P__260  (.L_HI(net260));
 sg13g2_tiehi \simon1.state[7]$_DFF_P__261  (.L_HI(net261));
 sg13g2_tiehi \simon1.tick_counter[0]$_SDFF_PP0__262  (.L_HI(net262));
 sg13g2_tiehi \simon1.tick_counter[10]$_SDFF_PP0__263  (.L_HI(net263));
 sg13g2_tiehi \simon1.tick_counter[11]$_SDFF_PP0__264  (.L_HI(net264));
 sg13g2_tiehi \simon1.tick_counter[12]$_SDFF_PP0__265  (.L_HI(net265));
 sg13g2_tiehi \simon1.tick_counter[13]$_SDFF_PP0__266  (.L_HI(net266));
 sg13g2_tiehi \simon1.tick_counter[14]$_SDFF_PP0__267  (.L_HI(net267));
 sg13g2_tiehi \simon1.tick_counter[15]$_SDFF_PP0__268  (.L_HI(net268));
 sg13g2_tiehi \simon1.tick_counter[1]$_SDFF_PP0__269  (.L_HI(net269));
 sg13g2_tiehi \simon1.tick_counter[2]$_SDFF_PP0__270  (.L_HI(net270));
 sg13g2_tiehi \simon1.tick_counter[3]$_SDFF_PP0__271  (.L_HI(net271));
 sg13g2_tiehi \simon1.tick_counter[4]$_SDFF_PP0__272  (.L_HI(net272));
 sg13g2_tiehi \simon1.tick_counter[5]$_SDFF_PP0__273  (.L_HI(net273));
 sg13g2_tiehi \simon1.tick_counter[6]$_SDFF_PP0__274  (.L_HI(net274));
 sg13g2_tiehi \simon1.tick_counter[7]$_SDFF_PP0__275  (.L_HI(net275));
 sg13g2_tiehi \simon1.tick_counter[8]$_SDFF_PP0__276  (.L_HI(net276));
 sg13g2_tiehi \simon1.tick_counter[9]$_SDFF_PP0__277  (.L_HI(net277));
 sg13g2_tiehi \simon1.tone_sequence_counter[0]$_DFFE_PP__278  (.L_HI(net278));
 sg13g2_tiehi \simon1.tone_sequence_counter[1]$_DFFE_PP__279  (.L_HI(net279));
 sg13g2_tiehi \simon1.tone_sequence_counter[2]$_DFFE_PP__280  (.L_HI(net280));
 sg13g2_tiehi \simon1.user_input[0]$_DFFE_PP__281  (.L_HI(net281));
 sg13g2_tiehi \simon1.user_input[1]$_DFFE_PP__282  (.L_HI(net282));
 sg13g2_tiehi \uio_out[0]$_DFF_P__283  (.L_HI(net283));
 sg13g2_tiehi \uio_out[1]$_DFF_P__284  (.L_HI(net284));
 sg13g2_tiehi \uio_out[2]$_DFF_P__285  (.L_HI(net285));
 sg13g2_tiehi \uio_out[3]$_DFF_P__286  (.L_HI(net286));
 sg13g2_tiehi \uio_out[4]$_DFF_P__287  (.L_HI(net287));
 sg13g2_tiehi \uio_out[5]$_DFF_P__288  (.L_HI(net288));
 sg13g2_tiehi \uio_out[6]$_DFF_P__289  (.L_HI(net289));
 sg13g2_tiehi \uo_out[0]$_SDFFE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \uo_out[1]$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \uo_out[2]$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_tiehi \uo_out[3]$_SDFFE_PN0P__293  (.L_HI(net293));
 sg13g2_tiehi \uo_out[5]$_DFF_P__294  (.L_HI(net294));
 sg13g2_tiehi \uo_out[6]$_DFF_P__295  (.L_HI(net295));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_inv_8 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_inv_8 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_inv_8 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_8 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_4_9_0_clk));
 sg13g2_buf_16 clkload10 (.A(clknet_4_10_0_clk));
 sg13g2_inv_8 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_8 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_inv_8 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_buf_16 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0109_));
 sg13g2_antennanp ANTENNA_2 (.A(_0109_));
 sg13g2_antennanp ANTENNA_3 (.A(_0111_));
 sg13g2_antennanp ANTENNA_4 (.A(_0111_));
 sg13g2_antennanp ANTENNA_5 (.A(_0112_));
 sg13g2_antennanp ANTENNA_6 (.A(_0112_));
 sg13g2_decap_8 FILLER_0_0_0 ();
 sg13g2_decap_8 FILLER_0_0_7 ();
 sg13g2_decap_8 FILLER_0_0_14 ();
 sg13g2_decap_8 FILLER_0_0_21 ();
 sg13g2_decap_8 FILLER_0_0_28 ();
 sg13g2_decap_8 FILLER_0_0_35 ();
 sg13g2_decap_8 FILLER_0_0_42 ();
 sg13g2_decap_8 FILLER_0_0_49 ();
 sg13g2_decap_8 FILLER_0_0_56 ();
 sg13g2_decap_8 FILLER_0_0_63 ();
 sg13g2_decap_8 FILLER_0_0_70 ();
 sg13g2_fill_2 FILLER_0_0_77 ();
 sg13g2_fill_2 FILLER_0_0_87 ();
 sg13g2_fill_2 FILLER_0_0_99 ();
 sg13g2_decap_4 FILLER_0_0_105 ();
 sg13g2_fill_1 FILLER_0_0_109 ();
 sg13g2_decap_8 FILLER_0_0_140 ();
 sg13g2_decap_8 FILLER_0_0_173 ();
 sg13g2_decap_8 FILLER_0_0_180 ();
 sg13g2_decap_8 FILLER_0_0_187 ();
 sg13g2_decap_8 FILLER_0_0_194 ();
 sg13g2_decap_8 FILLER_0_0_201 ();
 sg13g2_decap_8 FILLER_0_0_208 ();
 sg13g2_decap_8 FILLER_0_0_215 ();
 sg13g2_decap_8 FILLER_0_0_222 ();
 sg13g2_decap_8 FILLER_0_0_229 ();
 sg13g2_decap_8 FILLER_0_0_236 ();
 sg13g2_decap_8 FILLER_0_0_243 ();
 sg13g2_decap_8 FILLER_0_0_250 ();
 sg13g2_decap_8 FILLER_0_0_257 ();
 sg13g2_decap_8 FILLER_0_0_264 ();
 sg13g2_decap_8 FILLER_0_0_271 ();
 sg13g2_decap_8 FILLER_0_0_278 ();
 sg13g2_decap_8 FILLER_0_0_285 ();
 sg13g2_decap_8 FILLER_0_0_292 ();
 sg13g2_decap_8 FILLER_0_0_299 ();
 sg13g2_decap_8 FILLER_0_0_306 ();
 sg13g2_decap_8 FILLER_0_0_313 ();
 sg13g2_fill_2 FILLER_0_0_320 ();
 sg13g2_fill_1 FILLER_0_0_322 ();
 sg13g2_decap_8 FILLER_0_1_0 ();
 sg13g2_decap_8 FILLER_0_1_7 ();
 sg13g2_decap_8 FILLER_0_1_14 ();
 sg13g2_decap_8 FILLER_0_1_21 ();
 sg13g2_decap_8 FILLER_0_1_28 ();
 sg13g2_decap_8 FILLER_0_1_35 ();
 sg13g2_decap_8 FILLER_0_1_42 ();
 sg13g2_decap_8 FILLER_0_1_49 ();
 sg13g2_decap_4 FILLER_0_1_56 ();
 sg13g2_fill_1 FILLER_0_1_104 ();
 sg13g2_decap_4 FILLER_0_1_151 ();
 sg13g2_decap_8 FILLER_0_1_159 ();
 sg13g2_fill_2 FILLER_0_1_166 ();
 sg13g2_decap_8 FILLER_0_1_172 ();
 sg13g2_decap_8 FILLER_0_1_179 ();
 sg13g2_decap_8 FILLER_0_1_186 ();
 sg13g2_decap_8 FILLER_0_1_193 ();
 sg13g2_decap_8 FILLER_0_1_200 ();
 sg13g2_decap_8 FILLER_0_1_207 ();
 sg13g2_decap_8 FILLER_0_1_214 ();
 sg13g2_decap_8 FILLER_0_1_221 ();
 sg13g2_decap_8 FILLER_0_1_228 ();
 sg13g2_decap_8 FILLER_0_1_235 ();
 sg13g2_decap_8 FILLER_0_1_242 ();
 sg13g2_decap_8 FILLER_0_1_249 ();
 sg13g2_decap_8 FILLER_0_1_256 ();
 sg13g2_decap_8 FILLER_0_1_263 ();
 sg13g2_decap_8 FILLER_0_1_270 ();
 sg13g2_decap_8 FILLER_0_1_277 ();
 sg13g2_decap_8 FILLER_0_1_284 ();
 sg13g2_decap_8 FILLER_0_1_291 ();
 sg13g2_decap_8 FILLER_0_1_298 ();
 sg13g2_decap_8 FILLER_0_1_305 ();
 sg13g2_decap_8 FILLER_0_1_312 ();
 sg13g2_decap_4 FILLER_0_1_319 ();
 sg13g2_decap_8 FILLER_0_2_0 ();
 sg13g2_decap_8 FILLER_0_2_7 ();
 sg13g2_decap_8 FILLER_0_2_14 ();
 sg13g2_decap_8 FILLER_0_2_21 ();
 sg13g2_decap_8 FILLER_0_2_28 ();
 sg13g2_decap_8 FILLER_0_2_35 ();
 sg13g2_decap_8 FILLER_0_2_42 ();
 sg13g2_decap_8 FILLER_0_2_49 ();
 sg13g2_fill_1 FILLER_0_2_56 ();
 sg13g2_fill_1 FILLER_0_2_93 ();
 sg13g2_decap_8 FILLER_0_2_128 ();
 sg13g2_decap_8 FILLER_0_2_185 ();
 sg13g2_decap_8 FILLER_0_2_192 ();
 sg13g2_decap_8 FILLER_0_2_199 ();
 sg13g2_decap_8 FILLER_0_2_206 ();
 sg13g2_decap_8 FILLER_0_2_213 ();
 sg13g2_decap_8 FILLER_0_2_220 ();
 sg13g2_decap_8 FILLER_0_2_227 ();
 sg13g2_decap_8 FILLER_0_2_234 ();
 sg13g2_decap_8 FILLER_0_2_241 ();
 sg13g2_decap_8 FILLER_0_2_248 ();
 sg13g2_decap_8 FILLER_0_2_255 ();
 sg13g2_decap_8 FILLER_0_2_262 ();
 sg13g2_decap_8 FILLER_0_2_269 ();
 sg13g2_decap_8 FILLER_0_2_276 ();
 sg13g2_decap_8 FILLER_0_2_283 ();
 sg13g2_decap_8 FILLER_0_2_290 ();
 sg13g2_decap_8 FILLER_0_2_297 ();
 sg13g2_decap_8 FILLER_0_2_304 ();
 sg13g2_decap_8 FILLER_0_2_311 ();
 sg13g2_decap_4 FILLER_0_2_318 ();
 sg13g2_fill_1 FILLER_0_2_322 ();
 sg13g2_decap_8 FILLER_0_3_0 ();
 sg13g2_decap_8 FILLER_0_3_7 ();
 sg13g2_decap_8 FILLER_0_3_14 ();
 sg13g2_decap_8 FILLER_0_3_21 ();
 sg13g2_decap_8 FILLER_0_3_28 ();
 sg13g2_decap_8 FILLER_0_3_35 ();
 sg13g2_decap_8 FILLER_0_3_42 ();
 sg13g2_decap_4 FILLER_0_3_49 ();
 sg13g2_fill_2 FILLER_0_3_129 ();
 sg13g2_fill_1 FILLER_0_3_131 ();
 sg13g2_decap_8 FILLER_0_3_179 ();
 sg13g2_decap_8 FILLER_0_3_186 ();
 sg13g2_decap_8 FILLER_0_3_193 ();
 sg13g2_decap_8 FILLER_0_3_200 ();
 sg13g2_decap_8 FILLER_0_3_207 ();
 sg13g2_decap_8 FILLER_0_3_214 ();
 sg13g2_decap_8 FILLER_0_3_221 ();
 sg13g2_decap_8 FILLER_0_3_228 ();
 sg13g2_decap_8 FILLER_0_3_235 ();
 sg13g2_decap_8 FILLER_0_3_242 ();
 sg13g2_decap_8 FILLER_0_3_249 ();
 sg13g2_decap_8 FILLER_0_3_256 ();
 sg13g2_decap_8 FILLER_0_3_263 ();
 sg13g2_decap_8 FILLER_0_3_270 ();
 sg13g2_decap_8 FILLER_0_3_277 ();
 sg13g2_decap_8 FILLER_0_3_284 ();
 sg13g2_decap_8 FILLER_0_3_291 ();
 sg13g2_decap_8 FILLER_0_3_298 ();
 sg13g2_decap_8 FILLER_0_3_305 ();
 sg13g2_decap_8 FILLER_0_3_312 ();
 sg13g2_decap_4 FILLER_0_3_319 ();
 sg13g2_decap_8 FILLER_0_4_0 ();
 sg13g2_decap_8 FILLER_0_4_7 ();
 sg13g2_decap_8 FILLER_0_4_14 ();
 sg13g2_decap_8 FILLER_0_4_21 ();
 sg13g2_decap_8 FILLER_0_4_28 ();
 sg13g2_decap_8 FILLER_0_4_35 ();
 sg13g2_fill_2 FILLER_0_4_42 ();
 sg13g2_fill_1 FILLER_0_4_80 ();
 sg13g2_fill_1 FILLER_0_4_86 ();
 sg13g2_fill_2 FILLER_0_4_96 ();
 sg13g2_fill_1 FILLER_0_4_98 ();
 sg13g2_decap_8 FILLER_0_4_183 ();
 sg13g2_decap_8 FILLER_0_4_190 ();
 sg13g2_decap_8 FILLER_0_4_197 ();
 sg13g2_decap_8 FILLER_0_4_204 ();
 sg13g2_decap_8 FILLER_0_4_211 ();
 sg13g2_decap_8 FILLER_0_4_218 ();
 sg13g2_decap_8 FILLER_0_4_225 ();
 sg13g2_decap_8 FILLER_0_4_232 ();
 sg13g2_decap_8 FILLER_0_4_239 ();
 sg13g2_decap_8 FILLER_0_4_246 ();
 sg13g2_decap_8 FILLER_0_4_253 ();
 sg13g2_decap_8 FILLER_0_4_260 ();
 sg13g2_decap_8 FILLER_0_4_267 ();
 sg13g2_decap_8 FILLER_0_4_274 ();
 sg13g2_decap_8 FILLER_0_4_281 ();
 sg13g2_decap_8 FILLER_0_4_288 ();
 sg13g2_decap_8 FILLER_0_4_295 ();
 sg13g2_decap_8 FILLER_0_4_302 ();
 sg13g2_decap_8 FILLER_0_4_309 ();
 sg13g2_decap_8 FILLER_0_4_316 ();
 sg13g2_decap_8 FILLER_0_5_0 ();
 sg13g2_decap_8 FILLER_0_5_7 ();
 sg13g2_decap_8 FILLER_0_5_14 ();
 sg13g2_decap_8 FILLER_0_5_21 ();
 sg13g2_decap_8 FILLER_0_5_28 ();
 sg13g2_fill_2 FILLER_0_5_35 ();
 sg13g2_fill_1 FILLER_0_5_98 ();
 sg13g2_decap_8 FILLER_0_5_175 ();
 sg13g2_decap_8 FILLER_0_5_182 ();
 sg13g2_decap_8 FILLER_0_5_189 ();
 sg13g2_decap_8 FILLER_0_5_196 ();
 sg13g2_decap_8 FILLER_0_5_203 ();
 sg13g2_decap_8 FILLER_0_5_210 ();
 sg13g2_decap_8 FILLER_0_5_217 ();
 sg13g2_decap_8 FILLER_0_5_224 ();
 sg13g2_decap_8 FILLER_0_5_231 ();
 sg13g2_decap_8 FILLER_0_5_238 ();
 sg13g2_decap_8 FILLER_0_5_245 ();
 sg13g2_decap_8 FILLER_0_5_252 ();
 sg13g2_decap_8 FILLER_0_5_259 ();
 sg13g2_decap_8 FILLER_0_5_266 ();
 sg13g2_decap_8 FILLER_0_5_273 ();
 sg13g2_decap_8 FILLER_0_5_280 ();
 sg13g2_decap_8 FILLER_0_5_287 ();
 sg13g2_decap_8 FILLER_0_5_294 ();
 sg13g2_decap_8 FILLER_0_5_301 ();
 sg13g2_decap_8 FILLER_0_5_308 ();
 sg13g2_decap_8 FILLER_0_5_315 ();
 sg13g2_fill_1 FILLER_0_5_322 ();
 sg13g2_decap_8 FILLER_0_6_0 ();
 sg13g2_decap_8 FILLER_0_6_7 ();
 sg13g2_decap_8 FILLER_0_6_14 ();
 sg13g2_decap_8 FILLER_0_6_21 ();
 sg13g2_decap_8 FILLER_0_6_28 ();
 sg13g2_decap_8 FILLER_0_6_35 ();
 sg13g2_fill_2 FILLER_0_6_42 ();
 sg13g2_fill_1 FILLER_0_6_44 ();
 sg13g2_fill_2 FILLER_0_6_75 ();
 sg13g2_fill_2 FILLER_0_6_173 ();
 sg13g2_decap_8 FILLER_0_6_179 ();
 sg13g2_decap_8 FILLER_0_6_186 ();
 sg13g2_decap_8 FILLER_0_6_193 ();
 sg13g2_decap_8 FILLER_0_6_200 ();
 sg13g2_decap_8 FILLER_0_6_207 ();
 sg13g2_decap_8 FILLER_0_6_214 ();
 sg13g2_decap_8 FILLER_0_6_221 ();
 sg13g2_decap_8 FILLER_0_6_228 ();
 sg13g2_decap_8 FILLER_0_6_235 ();
 sg13g2_decap_8 FILLER_0_6_242 ();
 sg13g2_decap_8 FILLER_0_6_249 ();
 sg13g2_decap_8 FILLER_0_6_256 ();
 sg13g2_decap_8 FILLER_0_6_263 ();
 sg13g2_decap_8 FILLER_0_6_270 ();
 sg13g2_decap_8 FILLER_0_6_277 ();
 sg13g2_decap_8 FILLER_0_6_284 ();
 sg13g2_decap_8 FILLER_0_6_291 ();
 sg13g2_decap_8 FILLER_0_6_298 ();
 sg13g2_decap_8 FILLER_0_6_305 ();
 sg13g2_decap_8 FILLER_0_6_312 ();
 sg13g2_decap_4 FILLER_0_6_319 ();
 sg13g2_decap_8 FILLER_0_7_0 ();
 sg13g2_decap_8 FILLER_0_7_7 ();
 sg13g2_decap_8 FILLER_0_7_14 ();
 sg13g2_decap_8 FILLER_0_7_21 ();
 sg13g2_decap_8 FILLER_0_7_28 ();
 sg13g2_fill_2 FILLER_0_7_75 ();
 sg13g2_fill_1 FILLER_0_7_77 ();
 sg13g2_fill_2 FILLER_0_7_162 ();
 sg13g2_decap_8 FILLER_0_7_190 ();
 sg13g2_decap_8 FILLER_0_7_197 ();
 sg13g2_decap_8 FILLER_0_7_204 ();
 sg13g2_decap_8 FILLER_0_7_211 ();
 sg13g2_decap_8 FILLER_0_7_218 ();
 sg13g2_decap_8 FILLER_0_7_225 ();
 sg13g2_decap_8 FILLER_0_7_232 ();
 sg13g2_decap_8 FILLER_0_7_239 ();
 sg13g2_decap_8 FILLER_0_7_246 ();
 sg13g2_decap_8 FILLER_0_7_253 ();
 sg13g2_decap_8 FILLER_0_7_260 ();
 sg13g2_decap_8 FILLER_0_7_267 ();
 sg13g2_decap_8 FILLER_0_7_274 ();
 sg13g2_decap_8 FILLER_0_7_281 ();
 sg13g2_decap_8 FILLER_0_7_288 ();
 sg13g2_decap_8 FILLER_0_7_295 ();
 sg13g2_decap_8 FILLER_0_7_302 ();
 sg13g2_decap_8 FILLER_0_7_309 ();
 sg13g2_decap_8 FILLER_0_7_316 ();
 sg13g2_decap_8 FILLER_0_8_0 ();
 sg13g2_decap_8 FILLER_0_8_7 ();
 sg13g2_decap_8 FILLER_0_8_14 ();
 sg13g2_decap_8 FILLER_0_8_21 ();
 sg13g2_decap_8 FILLER_0_8_28 ();
 sg13g2_decap_4 FILLER_0_8_35 ();
 sg13g2_fill_1 FILLER_0_8_39 ();
 sg13g2_fill_1 FILLER_0_8_83 ();
 sg13g2_fill_1 FILLER_0_8_114 ();
 sg13g2_fill_2 FILLER_0_8_125 ();
 sg13g2_fill_2 FILLER_0_8_163 ();
 sg13g2_decap_8 FILLER_0_8_195 ();
 sg13g2_decap_8 FILLER_0_8_202 ();
 sg13g2_decap_8 FILLER_0_8_209 ();
 sg13g2_decap_8 FILLER_0_8_216 ();
 sg13g2_decap_8 FILLER_0_8_223 ();
 sg13g2_decap_8 FILLER_0_8_230 ();
 sg13g2_decap_8 FILLER_0_8_237 ();
 sg13g2_decap_8 FILLER_0_8_244 ();
 sg13g2_decap_8 FILLER_0_8_251 ();
 sg13g2_decap_8 FILLER_0_8_258 ();
 sg13g2_decap_8 FILLER_0_8_265 ();
 sg13g2_decap_8 FILLER_0_8_272 ();
 sg13g2_decap_8 FILLER_0_8_279 ();
 sg13g2_decap_8 FILLER_0_8_286 ();
 sg13g2_decap_8 FILLER_0_8_293 ();
 sg13g2_decap_8 FILLER_0_8_300 ();
 sg13g2_decap_8 FILLER_0_8_307 ();
 sg13g2_decap_8 FILLER_0_8_314 ();
 sg13g2_fill_2 FILLER_0_8_321 ();
 sg13g2_decap_8 FILLER_0_9_0 ();
 sg13g2_decap_8 FILLER_0_9_7 ();
 sg13g2_decap_8 FILLER_0_9_14 ();
 sg13g2_decap_8 FILLER_0_9_21 ();
 sg13g2_decap_8 FILLER_0_9_28 ();
 sg13g2_fill_2 FILLER_0_9_35 ();
 sg13g2_fill_1 FILLER_0_9_37 ();
 sg13g2_fill_2 FILLER_0_9_74 ();
 sg13g2_fill_1 FILLER_0_9_76 ();
 sg13g2_fill_1 FILLER_0_9_147 ();
 sg13g2_fill_2 FILLER_0_9_162 ();
 sg13g2_decap_8 FILLER_0_9_190 ();
 sg13g2_decap_8 FILLER_0_9_197 ();
 sg13g2_decap_8 FILLER_0_9_204 ();
 sg13g2_decap_8 FILLER_0_9_211 ();
 sg13g2_decap_8 FILLER_0_9_218 ();
 sg13g2_decap_8 FILLER_0_9_225 ();
 sg13g2_decap_8 FILLER_0_9_232 ();
 sg13g2_decap_8 FILLER_0_9_239 ();
 sg13g2_decap_8 FILLER_0_9_246 ();
 sg13g2_decap_8 FILLER_0_9_253 ();
 sg13g2_decap_8 FILLER_0_9_260 ();
 sg13g2_decap_8 FILLER_0_9_267 ();
 sg13g2_decap_8 FILLER_0_9_274 ();
 sg13g2_decap_8 FILLER_0_9_281 ();
 sg13g2_decap_8 FILLER_0_9_288 ();
 sg13g2_decap_8 FILLER_0_9_295 ();
 sg13g2_decap_8 FILLER_0_9_302 ();
 sg13g2_decap_8 FILLER_0_9_309 ();
 sg13g2_decap_8 FILLER_0_9_316 ();
 sg13g2_decap_8 FILLER_0_10_0 ();
 sg13g2_decap_8 FILLER_0_10_7 ();
 sg13g2_decap_8 FILLER_0_10_14 ();
 sg13g2_decap_8 FILLER_0_10_21 ();
 sg13g2_decap_8 FILLER_0_10_28 ();
 sg13g2_fill_1 FILLER_0_10_168 ();
 sg13g2_fill_1 FILLER_0_10_173 ();
 sg13g2_fill_1 FILLER_0_10_200 ();
 sg13g2_decap_8 FILLER_0_10_205 ();
 sg13g2_decap_8 FILLER_0_10_212 ();
 sg13g2_decap_8 FILLER_0_10_219 ();
 sg13g2_decap_8 FILLER_0_10_226 ();
 sg13g2_decap_8 FILLER_0_10_233 ();
 sg13g2_decap_8 FILLER_0_10_240 ();
 sg13g2_decap_8 FILLER_0_10_247 ();
 sg13g2_decap_8 FILLER_0_10_254 ();
 sg13g2_decap_8 FILLER_0_10_261 ();
 sg13g2_decap_8 FILLER_0_10_268 ();
 sg13g2_decap_8 FILLER_0_10_275 ();
 sg13g2_decap_8 FILLER_0_10_282 ();
 sg13g2_decap_8 FILLER_0_10_289 ();
 sg13g2_decap_8 FILLER_0_10_296 ();
 sg13g2_decap_8 FILLER_0_10_303 ();
 sg13g2_decap_8 FILLER_0_10_310 ();
 sg13g2_decap_4 FILLER_0_10_317 ();
 sg13g2_fill_2 FILLER_0_10_321 ();
 sg13g2_decap_8 FILLER_0_11_0 ();
 sg13g2_decap_8 FILLER_0_11_7 ();
 sg13g2_decap_8 FILLER_0_11_14 ();
 sg13g2_decap_8 FILLER_0_11_21 ();
 sg13g2_fill_2 FILLER_0_11_28 ();
 sg13g2_fill_2 FILLER_0_11_38 ();
 sg13g2_fill_1 FILLER_0_11_101 ();
 sg13g2_decap_4 FILLER_0_11_171 ();
 sg13g2_fill_1 FILLER_0_11_175 ();
 sg13g2_decap_4 FILLER_0_11_189 ();
 sg13g2_fill_1 FILLER_0_11_193 ();
 sg13g2_decap_8 FILLER_0_11_220 ();
 sg13g2_decap_8 FILLER_0_11_227 ();
 sg13g2_decap_8 FILLER_0_11_234 ();
 sg13g2_decap_8 FILLER_0_11_241 ();
 sg13g2_decap_8 FILLER_0_11_248 ();
 sg13g2_decap_8 FILLER_0_11_255 ();
 sg13g2_decap_8 FILLER_0_11_262 ();
 sg13g2_decap_8 FILLER_0_11_269 ();
 sg13g2_decap_8 FILLER_0_11_276 ();
 sg13g2_decap_8 FILLER_0_11_283 ();
 sg13g2_decap_8 FILLER_0_11_290 ();
 sg13g2_decap_8 FILLER_0_11_297 ();
 sg13g2_decap_8 FILLER_0_11_304 ();
 sg13g2_decap_8 FILLER_0_11_311 ();
 sg13g2_decap_4 FILLER_0_11_318 ();
 sg13g2_fill_1 FILLER_0_11_322 ();
 sg13g2_decap_8 FILLER_0_12_0 ();
 sg13g2_decap_8 FILLER_0_12_7 ();
 sg13g2_decap_8 FILLER_0_12_14 ();
 sg13g2_decap_8 FILLER_0_12_21 ();
 sg13g2_fill_2 FILLER_0_12_28 ();
 sg13g2_fill_2 FILLER_0_12_95 ();
 sg13g2_fill_1 FILLER_0_12_141 ();
 sg13g2_fill_2 FILLER_0_12_147 ();
 sg13g2_decap_8 FILLER_0_12_195 ();
 sg13g2_decap_8 FILLER_0_12_202 ();
 sg13g2_decap_8 FILLER_0_12_209 ();
 sg13g2_decap_8 FILLER_0_12_216 ();
 sg13g2_decap_8 FILLER_0_12_223 ();
 sg13g2_decap_8 FILLER_0_12_230 ();
 sg13g2_decap_8 FILLER_0_12_237 ();
 sg13g2_decap_8 FILLER_0_12_244 ();
 sg13g2_decap_8 FILLER_0_12_251 ();
 sg13g2_decap_8 FILLER_0_12_258 ();
 sg13g2_decap_8 FILLER_0_12_265 ();
 sg13g2_decap_8 FILLER_0_12_272 ();
 sg13g2_decap_8 FILLER_0_12_279 ();
 sg13g2_decap_8 FILLER_0_12_286 ();
 sg13g2_decap_8 FILLER_0_12_293 ();
 sg13g2_decap_8 FILLER_0_12_300 ();
 sg13g2_decap_8 FILLER_0_12_307 ();
 sg13g2_decap_8 FILLER_0_12_314 ();
 sg13g2_fill_2 FILLER_0_12_321 ();
 sg13g2_decap_8 FILLER_0_13_0 ();
 sg13g2_decap_8 FILLER_0_13_7 ();
 sg13g2_decap_8 FILLER_0_13_14 ();
 sg13g2_decap_4 FILLER_0_13_21 ();
 sg13g2_fill_2 FILLER_0_13_25 ();
 sg13g2_decap_4 FILLER_0_13_31 ();
 sg13g2_fill_1 FILLER_0_13_35 ();
 sg13g2_fill_1 FILLER_0_13_108 ();
 sg13g2_fill_2 FILLER_0_13_143 ();
 sg13g2_decap_8 FILLER_0_13_185 ();
 sg13g2_decap_8 FILLER_0_13_192 ();
 sg13g2_decap_8 FILLER_0_13_199 ();
 sg13g2_decap_8 FILLER_0_13_206 ();
 sg13g2_decap_8 FILLER_0_13_213 ();
 sg13g2_decap_8 FILLER_0_13_220 ();
 sg13g2_decap_8 FILLER_0_13_227 ();
 sg13g2_decap_8 FILLER_0_13_234 ();
 sg13g2_decap_8 FILLER_0_13_241 ();
 sg13g2_decap_8 FILLER_0_13_248 ();
 sg13g2_decap_8 FILLER_0_13_255 ();
 sg13g2_decap_8 FILLER_0_13_262 ();
 sg13g2_decap_8 FILLER_0_13_269 ();
 sg13g2_decap_8 FILLER_0_13_276 ();
 sg13g2_decap_8 FILLER_0_13_283 ();
 sg13g2_decap_8 FILLER_0_13_290 ();
 sg13g2_decap_8 FILLER_0_13_297 ();
 sg13g2_decap_8 FILLER_0_13_304 ();
 sg13g2_decap_8 FILLER_0_13_311 ();
 sg13g2_decap_4 FILLER_0_13_318 ();
 sg13g2_fill_1 FILLER_0_13_322 ();
 sg13g2_decap_8 FILLER_0_14_0 ();
 sg13g2_decap_8 FILLER_0_14_7 ();
 sg13g2_decap_8 FILLER_0_14_14 ();
 sg13g2_decap_8 FILLER_0_14_21 ();
 sg13g2_decap_8 FILLER_0_14_28 ();
 sg13g2_fill_1 FILLER_0_14_35 ();
 sg13g2_decap_8 FILLER_0_14_189 ();
 sg13g2_decap_8 FILLER_0_14_196 ();
 sg13g2_decap_8 FILLER_0_14_203 ();
 sg13g2_decap_8 FILLER_0_14_210 ();
 sg13g2_decap_8 FILLER_0_14_217 ();
 sg13g2_decap_8 FILLER_0_14_224 ();
 sg13g2_decap_8 FILLER_0_14_231 ();
 sg13g2_decap_8 FILLER_0_14_238 ();
 sg13g2_decap_8 FILLER_0_14_245 ();
 sg13g2_decap_8 FILLER_0_14_252 ();
 sg13g2_decap_8 FILLER_0_14_259 ();
 sg13g2_decap_8 FILLER_0_14_266 ();
 sg13g2_decap_8 FILLER_0_14_273 ();
 sg13g2_decap_8 FILLER_0_14_280 ();
 sg13g2_decap_8 FILLER_0_14_287 ();
 sg13g2_decap_8 FILLER_0_14_294 ();
 sg13g2_decap_8 FILLER_0_14_301 ();
 sg13g2_decap_8 FILLER_0_14_308 ();
 sg13g2_decap_8 FILLER_0_14_315 ();
 sg13g2_fill_1 FILLER_0_14_322 ();
 sg13g2_decap_8 FILLER_0_15_0 ();
 sg13g2_decap_8 FILLER_0_15_7 ();
 sg13g2_decap_8 FILLER_0_15_14 ();
 sg13g2_decap_8 FILLER_0_15_21 ();
 sg13g2_decap_4 FILLER_0_15_28 ();
 sg13g2_fill_2 FILLER_0_15_106 ();
 sg13g2_fill_1 FILLER_0_15_118 ();
 sg13g2_decap_8 FILLER_0_15_189 ();
 sg13g2_decap_8 FILLER_0_15_196 ();
 sg13g2_decap_8 FILLER_0_15_203 ();
 sg13g2_decap_8 FILLER_0_15_210 ();
 sg13g2_decap_8 FILLER_0_15_217 ();
 sg13g2_decap_8 FILLER_0_15_224 ();
 sg13g2_decap_8 FILLER_0_15_231 ();
 sg13g2_decap_8 FILLER_0_15_238 ();
 sg13g2_decap_8 FILLER_0_15_245 ();
 sg13g2_decap_8 FILLER_0_15_252 ();
 sg13g2_decap_8 FILLER_0_15_259 ();
 sg13g2_decap_8 FILLER_0_15_266 ();
 sg13g2_decap_8 FILLER_0_15_273 ();
 sg13g2_decap_8 FILLER_0_15_280 ();
 sg13g2_decap_8 FILLER_0_15_287 ();
 sg13g2_decap_8 FILLER_0_15_294 ();
 sg13g2_decap_8 FILLER_0_15_301 ();
 sg13g2_decap_8 FILLER_0_15_308 ();
 sg13g2_decap_8 FILLER_0_15_315 ();
 sg13g2_fill_1 FILLER_0_15_322 ();
 sg13g2_decap_8 FILLER_0_16_0 ();
 sg13g2_decap_8 FILLER_0_16_7 ();
 sg13g2_decap_8 FILLER_0_16_14 ();
 sg13g2_decap_8 FILLER_0_16_21 ();
 sg13g2_decap_8 FILLER_0_16_28 ();
 sg13g2_decap_4 FILLER_0_16_35 ();
 sg13g2_fill_1 FILLER_0_16_39 ();
 sg13g2_fill_2 FILLER_0_16_97 ();
 sg13g2_fill_1 FILLER_0_16_138 ();
 sg13g2_fill_1 FILLER_0_16_170 ();
 sg13g2_fill_1 FILLER_0_16_175 ();
 sg13g2_decap_8 FILLER_0_16_202 ();
 sg13g2_decap_8 FILLER_0_16_209 ();
 sg13g2_decap_8 FILLER_0_16_216 ();
 sg13g2_decap_8 FILLER_0_16_223 ();
 sg13g2_decap_8 FILLER_0_16_230 ();
 sg13g2_decap_8 FILLER_0_16_237 ();
 sg13g2_decap_8 FILLER_0_16_244 ();
 sg13g2_decap_8 FILLER_0_16_251 ();
 sg13g2_decap_8 FILLER_0_16_258 ();
 sg13g2_decap_8 FILLER_0_16_265 ();
 sg13g2_decap_8 FILLER_0_16_272 ();
 sg13g2_decap_8 FILLER_0_16_279 ();
 sg13g2_decap_8 FILLER_0_16_286 ();
 sg13g2_decap_8 FILLER_0_16_293 ();
 sg13g2_decap_8 FILLER_0_16_300 ();
 sg13g2_decap_8 FILLER_0_16_307 ();
 sg13g2_decap_8 FILLER_0_16_314 ();
 sg13g2_fill_2 FILLER_0_16_321 ();
 sg13g2_decap_8 FILLER_0_17_0 ();
 sg13g2_decap_8 FILLER_0_17_7 ();
 sg13g2_decap_8 FILLER_0_17_14 ();
 sg13g2_decap_8 FILLER_0_17_21 ();
 sg13g2_decap_8 FILLER_0_17_28 ();
 sg13g2_decap_4 FILLER_0_17_35 ();
 sg13g2_fill_2 FILLER_0_17_116 ();
 sg13g2_fill_1 FILLER_0_17_148 ();
 sg13g2_decap_8 FILLER_0_17_159 ();
 sg13g2_decap_8 FILLER_0_17_166 ();
 sg13g2_decap_8 FILLER_0_17_173 ();
 sg13g2_decap_4 FILLER_0_17_180 ();
 sg13g2_decap_8 FILLER_0_17_188 ();
 sg13g2_decap_8 FILLER_0_17_195 ();
 sg13g2_decap_8 FILLER_0_17_202 ();
 sg13g2_decap_8 FILLER_0_17_209 ();
 sg13g2_decap_8 FILLER_0_17_216 ();
 sg13g2_decap_8 FILLER_0_17_223 ();
 sg13g2_decap_8 FILLER_0_17_230 ();
 sg13g2_decap_8 FILLER_0_17_237 ();
 sg13g2_decap_8 FILLER_0_17_244 ();
 sg13g2_decap_8 FILLER_0_17_251 ();
 sg13g2_decap_8 FILLER_0_17_258 ();
 sg13g2_decap_8 FILLER_0_17_265 ();
 sg13g2_decap_8 FILLER_0_17_272 ();
 sg13g2_decap_8 FILLER_0_17_279 ();
 sg13g2_decap_8 FILLER_0_17_286 ();
 sg13g2_decap_8 FILLER_0_17_293 ();
 sg13g2_decap_8 FILLER_0_17_300 ();
 sg13g2_decap_8 FILLER_0_17_307 ();
 sg13g2_decap_8 FILLER_0_17_314 ();
 sg13g2_fill_2 FILLER_0_17_321 ();
 sg13g2_decap_8 FILLER_0_18_0 ();
 sg13g2_decap_8 FILLER_0_18_7 ();
 sg13g2_decap_8 FILLER_0_18_14 ();
 sg13g2_decap_8 FILLER_0_18_21 ();
 sg13g2_decap_8 FILLER_0_18_28 ();
 sg13g2_decap_8 FILLER_0_18_35 ();
 sg13g2_fill_1 FILLER_0_18_68 ();
 sg13g2_fill_1 FILLER_0_18_84 ();
 sg13g2_fill_2 FILLER_0_18_113 ();
 sg13g2_decap_8 FILLER_0_18_182 ();
 sg13g2_decap_8 FILLER_0_18_189 ();
 sg13g2_decap_8 FILLER_0_18_196 ();
 sg13g2_decap_8 FILLER_0_18_203 ();
 sg13g2_decap_8 FILLER_0_18_210 ();
 sg13g2_decap_8 FILLER_0_18_217 ();
 sg13g2_decap_8 FILLER_0_18_224 ();
 sg13g2_decap_8 FILLER_0_18_231 ();
 sg13g2_decap_8 FILLER_0_18_238 ();
 sg13g2_decap_8 FILLER_0_18_245 ();
 sg13g2_decap_8 FILLER_0_18_252 ();
 sg13g2_decap_8 FILLER_0_18_259 ();
 sg13g2_decap_8 FILLER_0_18_266 ();
 sg13g2_decap_8 FILLER_0_18_273 ();
 sg13g2_decap_8 FILLER_0_18_280 ();
 sg13g2_decap_8 FILLER_0_18_287 ();
 sg13g2_decap_8 FILLER_0_18_294 ();
 sg13g2_decap_8 FILLER_0_18_301 ();
 sg13g2_decap_8 FILLER_0_18_308 ();
 sg13g2_decap_8 FILLER_0_18_315 ();
 sg13g2_fill_1 FILLER_0_18_322 ();
 sg13g2_decap_8 FILLER_0_19_0 ();
 sg13g2_decap_8 FILLER_0_19_7 ();
 sg13g2_fill_2 FILLER_0_19_14 ();
 sg13g2_decap_4 FILLER_0_19_42 ();
 sg13g2_fill_1 FILLER_0_19_46 ();
 sg13g2_fill_1 FILLER_0_19_51 ();
 sg13g2_fill_2 FILLER_0_19_62 ();
 sg13g2_fill_2 FILLER_0_19_78 ();
 sg13g2_fill_1 FILLER_0_19_80 ();
 sg13g2_fill_2 FILLER_0_19_91 ();
 sg13g2_fill_1 FILLER_0_19_93 ();
 sg13g2_fill_1 FILLER_0_19_135 ();
 sg13g2_fill_1 FILLER_0_19_157 ();
 sg13g2_decap_8 FILLER_0_19_184 ();
 sg13g2_decap_8 FILLER_0_19_191 ();
 sg13g2_decap_8 FILLER_0_19_198 ();
 sg13g2_decap_8 FILLER_0_19_205 ();
 sg13g2_decap_8 FILLER_0_19_212 ();
 sg13g2_decap_8 FILLER_0_19_219 ();
 sg13g2_decap_8 FILLER_0_19_226 ();
 sg13g2_decap_8 FILLER_0_19_233 ();
 sg13g2_decap_8 FILLER_0_19_240 ();
 sg13g2_decap_8 FILLER_0_19_247 ();
 sg13g2_decap_8 FILLER_0_19_254 ();
 sg13g2_decap_8 FILLER_0_19_261 ();
 sg13g2_decap_8 FILLER_0_19_268 ();
 sg13g2_decap_8 FILLER_0_19_275 ();
 sg13g2_decap_8 FILLER_0_19_282 ();
 sg13g2_decap_8 FILLER_0_19_289 ();
 sg13g2_decap_8 FILLER_0_19_296 ();
 sg13g2_decap_8 FILLER_0_19_303 ();
 sg13g2_decap_8 FILLER_0_19_310 ();
 sg13g2_decap_4 FILLER_0_19_317 ();
 sg13g2_fill_2 FILLER_0_19_321 ();
 sg13g2_decap_8 FILLER_0_20_0 ();
 sg13g2_decap_8 FILLER_0_20_7 ();
 sg13g2_decap_4 FILLER_0_20_14 ();
 sg13g2_fill_2 FILLER_0_20_18 ();
 sg13g2_decap_8 FILLER_0_20_24 ();
 sg13g2_fill_2 FILLER_0_20_51 ();
 sg13g2_fill_1 FILLER_0_20_53 ();
 sg13g2_fill_2 FILLER_0_20_101 ();
 sg13g2_fill_1 FILLER_0_20_103 ();
 sg13g2_fill_2 FILLER_0_20_114 ();
 sg13g2_fill_1 FILLER_0_20_142 ();
 sg13g2_decap_4 FILLER_0_20_172 ();
 sg13g2_fill_2 FILLER_0_20_176 ();
 sg13g2_decap_8 FILLER_0_20_183 ();
 sg13g2_decap_8 FILLER_0_20_190 ();
 sg13g2_decap_8 FILLER_0_20_197 ();
 sg13g2_decap_8 FILLER_0_20_204 ();
 sg13g2_decap_8 FILLER_0_20_211 ();
 sg13g2_decap_8 FILLER_0_20_218 ();
 sg13g2_decap_8 FILLER_0_20_225 ();
 sg13g2_decap_8 FILLER_0_20_232 ();
 sg13g2_decap_8 FILLER_0_20_239 ();
 sg13g2_decap_8 FILLER_0_20_246 ();
 sg13g2_decap_8 FILLER_0_20_253 ();
 sg13g2_decap_8 FILLER_0_20_260 ();
 sg13g2_decap_8 FILLER_0_20_267 ();
 sg13g2_decap_8 FILLER_0_20_274 ();
 sg13g2_fill_2 FILLER_0_20_285 ();
 sg13g2_fill_1 FILLER_0_20_287 ();
 sg13g2_fill_1 FILLER_0_20_292 ();
 sg13g2_decap_8 FILLER_0_21_0 ();
 sg13g2_decap_8 FILLER_0_21_7 ();
 sg13g2_decap_8 FILLER_0_21_14 ();
 sg13g2_decap_8 FILLER_0_21_21 ();
 sg13g2_decap_4 FILLER_0_21_28 ();
 sg13g2_fill_2 FILLER_0_21_32 ();
 sg13g2_fill_1 FILLER_0_21_64 ();
 sg13g2_fill_2 FILLER_0_21_92 ();
 sg13g2_fill_1 FILLER_0_21_94 ();
 sg13g2_fill_2 FILLER_0_21_142 ();
 sg13g2_fill_1 FILLER_0_21_165 ();
 sg13g2_decap_4 FILLER_0_21_174 ();
 sg13g2_decap_8 FILLER_0_21_188 ();
 sg13g2_decap_8 FILLER_0_21_195 ();
 sg13g2_decap_8 FILLER_0_21_202 ();
 sg13g2_fill_2 FILLER_0_21_209 ();
 sg13g2_fill_1 FILLER_0_21_211 ();
 sg13g2_decap_8 FILLER_0_21_227 ();
 sg13g2_decap_8 FILLER_0_21_234 ();
 sg13g2_decap_8 FILLER_0_21_241 ();
 sg13g2_decap_8 FILLER_0_21_248 ();
 sg13g2_decap_8 FILLER_0_21_255 ();
 sg13g2_decap_4 FILLER_0_21_262 ();
 sg13g2_decap_4 FILLER_0_21_270 ();
 sg13g2_fill_2 FILLER_0_21_312 ();
 sg13g2_fill_1 FILLER_0_21_314 ();
 sg13g2_decap_8 FILLER_0_22_0 ();
 sg13g2_decap_8 FILLER_0_22_7 ();
 sg13g2_decap_8 FILLER_0_22_14 ();
 sg13g2_decap_8 FILLER_0_22_21 ();
 sg13g2_decap_8 FILLER_0_22_28 ();
 sg13g2_fill_2 FILLER_0_22_35 ();
 sg13g2_fill_1 FILLER_0_22_37 ();
 sg13g2_decap_8 FILLER_0_22_181 ();
 sg13g2_decap_8 FILLER_0_22_188 ();
 sg13g2_decap_8 FILLER_0_22_195 ();
 sg13g2_decap_8 FILLER_0_22_202 ();
 sg13g2_decap_8 FILLER_0_22_209 ();
 sg13g2_decap_8 FILLER_0_22_216 ();
 sg13g2_decap_8 FILLER_0_22_223 ();
 sg13g2_decap_8 FILLER_0_22_230 ();
 sg13g2_decap_8 FILLER_0_22_237 ();
 sg13g2_decap_8 FILLER_0_22_244 ();
 sg13g2_decap_8 FILLER_0_22_251 ();
 sg13g2_fill_1 FILLER_0_22_258 ();
 sg13g2_fill_1 FILLER_0_22_307 ();
 sg13g2_fill_2 FILLER_0_22_315 ();
 sg13g2_fill_1 FILLER_0_22_317 ();
 sg13g2_fill_1 FILLER_0_22_322 ();
 sg13g2_decap_8 FILLER_0_23_0 ();
 sg13g2_decap_8 FILLER_0_23_7 ();
 sg13g2_decap_8 FILLER_0_23_14 ();
 sg13g2_decap_8 FILLER_0_23_21 ();
 sg13g2_decap_4 FILLER_0_23_28 ();
 sg13g2_fill_1 FILLER_0_23_32 ();
 sg13g2_fill_1 FILLER_0_23_100 ();
 sg13g2_fill_1 FILLER_0_23_113 ();
 sg13g2_fill_1 FILLER_0_23_140 ();
 sg13g2_fill_2 FILLER_0_23_177 ();
 sg13g2_decap_8 FILLER_0_23_183 ();
 sg13g2_decap_8 FILLER_0_23_190 ();
 sg13g2_decap_8 FILLER_0_23_197 ();
 sg13g2_decap_8 FILLER_0_23_204 ();
 sg13g2_decap_8 FILLER_0_23_211 ();
 sg13g2_decap_8 FILLER_0_23_218 ();
 sg13g2_decap_8 FILLER_0_23_225 ();
 sg13g2_decap_8 FILLER_0_23_232 ();
 sg13g2_decap_8 FILLER_0_23_239 ();
 sg13g2_decap_8 FILLER_0_23_246 ();
 sg13g2_decap_4 FILLER_0_23_253 ();
 sg13g2_fill_2 FILLER_0_23_257 ();
 sg13g2_fill_2 FILLER_0_23_295 ();
 sg13g2_decap_8 FILLER_0_24_0 ();
 sg13g2_decap_8 FILLER_0_24_7 ();
 sg13g2_decap_8 FILLER_0_24_14 ();
 sg13g2_decap_8 FILLER_0_24_21 ();
 sg13g2_decap_4 FILLER_0_24_28 ();
 sg13g2_fill_1 FILLER_0_24_32 ();
 sg13g2_fill_2 FILLER_0_24_78 ();
 sg13g2_fill_1 FILLER_0_24_80 ();
 sg13g2_fill_1 FILLER_0_24_109 ();
 sg13g2_fill_1 FILLER_0_24_114 ();
 sg13g2_decap_8 FILLER_0_24_181 ();
 sg13g2_decap_8 FILLER_0_24_188 ();
 sg13g2_decap_8 FILLER_0_24_195 ();
 sg13g2_decap_8 FILLER_0_24_202 ();
 sg13g2_decap_8 FILLER_0_24_209 ();
 sg13g2_decap_8 FILLER_0_24_216 ();
 sg13g2_decap_8 FILLER_0_24_223 ();
 sg13g2_decap_8 FILLER_0_24_230 ();
 sg13g2_decap_4 FILLER_0_24_237 ();
 sg13g2_fill_1 FILLER_0_24_258 ();
 sg13g2_fill_2 FILLER_0_24_294 ();
 sg13g2_fill_1 FILLER_0_24_296 ();
 sg13g2_decap_8 FILLER_0_25_0 ();
 sg13g2_decap_8 FILLER_0_25_7 ();
 sg13g2_decap_8 FILLER_0_25_14 ();
 sg13g2_decap_8 FILLER_0_25_21 ();
 sg13g2_decap_8 FILLER_0_25_28 ();
 sg13g2_decap_8 FILLER_0_25_35 ();
 sg13g2_decap_4 FILLER_0_25_42 ();
 sg13g2_fill_1 FILLER_0_25_46 ();
 sg13g2_fill_1 FILLER_0_25_94 ();
 sg13g2_fill_1 FILLER_0_25_100 ();
 sg13g2_fill_1 FILLER_0_25_106 ();
 sg13g2_fill_2 FILLER_0_25_111 ();
 sg13g2_fill_1 FILLER_0_25_139 ();
 sg13g2_decap_8 FILLER_0_25_170 ();
 sg13g2_decap_8 FILLER_0_25_177 ();
 sg13g2_decap_8 FILLER_0_25_184 ();
 sg13g2_decap_8 FILLER_0_25_191 ();
 sg13g2_decap_8 FILLER_0_25_198 ();
 sg13g2_decap_8 FILLER_0_25_205 ();
 sg13g2_fill_2 FILLER_0_25_212 ();
 sg13g2_decap_8 FILLER_0_25_217 ();
 sg13g2_decap_8 FILLER_0_25_224 ();
 sg13g2_decap_8 FILLER_0_25_231 ();
 sg13g2_fill_2 FILLER_0_25_238 ();
 sg13g2_fill_2 FILLER_0_25_271 ();
 sg13g2_fill_1 FILLER_0_25_273 ();
 sg13g2_fill_1 FILLER_0_25_295 ();
 sg13g2_fill_2 FILLER_0_25_321 ();
 sg13g2_decap_8 FILLER_0_26_0 ();
 sg13g2_decap_8 FILLER_0_26_7 ();
 sg13g2_decap_8 FILLER_0_26_14 ();
 sg13g2_decap_8 FILLER_0_26_21 ();
 sg13g2_decap_8 FILLER_0_26_28 ();
 sg13g2_decap_8 FILLER_0_26_35 ();
 sg13g2_fill_2 FILLER_0_26_42 ();
 sg13g2_fill_1 FILLER_0_26_44 ();
 sg13g2_decap_8 FILLER_0_26_49 ();
 sg13g2_fill_2 FILLER_0_26_56 ();
 sg13g2_fill_1 FILLER_0_26_58 ();
 sg13g2_fill_1 FILLER_0_26_125 ();
 sg13g2_fill_2 FILLER_0_26_138 ();
 sg13g2_decap_8 FILLER_0_26_170 ();
 sg13g2_decap_8 FILLER_0_26_177 ();
 sg13g2_decap_8 FILLER_0_26_184 ();
 sg13g2_decap_8 FILLER_0_26_191 ();
 sg13g2_decap_8 FILLER_0_26_198 ();
 sg13g2_decap_8 FILLER_0_26_205 ();
 sg13g2_decap_8 FILLER_0_26_212 ();
 sg13g2_decap_8 FILLER_0_26_219 ();
 sg13g2_decap_8 FILLER_0_26_226 ();
 sg13g2_decap_4 FILLER_0_26_233 ();
 sg13g2_fill_2 FILLER_0_26_259 ();
 sg13g2_fill_1 FILLER_0_26_266 ();
 sg13g2_decap_8 FILLER_0_27_0 ();
 sg13g2_decap_8 FILLER_0_27_7 ();
 sg13g2_decap_8 FILLER_0_27_14 ();
 sg13g2_decap_8 FILLER_0_27_21 ();
 sg13g2_decap_8 FILLER_0_27_28 ();
 sg13g2_fill_2 FILLER_0_27_35 ();
 sg13g2_fill_1 FILLER_0_27_37 ();
 sg13g2_decap_4 FILLER_0_27_64 ();
 sg13g2_fill_2 FILLER_0_27_68 ();
 sg13g2_fill_1 FILLER_0_27_101 ();
 sg13g2_fill_2 FILLER_0_27_136 ();
 sg13g2_decap_8 FILLER_0_27_164 ();
 sg13g2_decap_8 FILLER_0_27_171 ();
 sg13g2_decap_8 FILLER_0_27_178 ();
 sg13g2_decap_8 FILLER_0_27_185 ();
 sg13g2_decap_8 FILLER_0_27_192 ();
 sg13g2_decap_8 FILLER_0_27_199 ();
 sg13g2_decap_8 FILLER_0_27_206 ();
 sg13g2_decap_8 FILLER_0_27_213 ();
 sg13g2_decap_8 FILLER_0_27_220 ();
 sg13g2_decap_8 FILLER_0_27_227 ();
 sg13g2_decap_8 FILLER_0_27_234 ();
 sg13g2_fill_1 FILLER_0_27_250 ();
 sg13g2_fill_1 FILLER_0_27_259 ();
 sg13g2_fill_2 FILLER_0_27_282 ();
 sg13g2_fill_1 FILLER_0_27_284 ();
 sg13g2_fill_1 FILLER_0_27_297 ();
 sg13g2_fill_1 FILLER_0_27_304 ();
 sg13g2_fill_1 FILLER_0_27_316 ();
 sg13g2_fill_1 FILLER_0_27_322 ();
 sg13g2_decap_8 FILLER_0_28_0 ();
 sg13g2_decap_8 FILLER_0_28_7 ();
 sg13g2_decap_8 FILLER_0_28_14 ();
 sg13g2_decap_4 FILLER_0_28_21 ();
 sg13g2_fill_2 FILLER_0_28_25 ();
 sg13g2_fill_1 FILLER_0_28_109 ();
 sg13g2_fill_1 FILLER_0_28_115 ();
 sg13g2_fill_2 FILLER_0_28_124 ();
 sg13g2_fill_2 FILLER_0_28_131 ();
 sg13g2_fill_2 FILLER_0_28_138 ();
 sg13g2_decap_8 FILLER_0_28_166 ();
 sg13g2_decap_8 FILLER_0_28_173 ();
 sg13g2_decap_8 FILLER_0_28_180 ();
 sg13g2_decap_8 FILLER_0_28_187 ();
 sg13g2_decap_8 FILLER_0_28_194 ();
 sg13g2_decap_8 FILLER_0_28_201 ();
 sg13g2_decap_8 FILLER_0_28_208 ();
 sg13g2_decap_8 FILLER_0_28_215 ();
 sg13g2_fill_1 FILLER_0_28_222 ();
 sg13g2_fill_2 FILLER_0_28_283 ();
 sg13g2_fill_2 FILLER_0_28_300 ();
 sg13g2_fill_1 FILLER_0_28_322 ();
 sg13g2_decap_8 FILLER_0_29_0 ();
 sg13g2_decap_8 FILLER_0_29_7 ();
 sg13g2_decap_8 FILLER_0_29_14 ();
 sg13g2_decap_8 FILLER_0_29_21 ();
 sg13g2_fill_2 FILLER_0_29_28 ();
 sg13g2_decap_4 FILLER_0_29_34 ();
 sg13g2_fill_1 FILLER_0_29_42 ();
 sg13g2_fill_1 FILLER_0_29_132 ();
 sg13g2_fill_1 FILLER_0_29_138 ();
 sg13g2_fill_2 FILLER_0_29_152 ();
 sg13g2_fill_1 FILLER_0_29_154 ();
 sg13g2_decap_8 FILLER_0_29_159 ();
 sg13g2_fill_2 FILLER_0_29_166 ();
 sg13g2_fill_1 FILLER_0_29_168 ();
 sg13g2_decap_8 FILLER_0_29_173 ();
 sg13g2_decap_8 FILLER_0_29_180 ();
 sg13g2_decap_8 FILLER_0_29_187 ();
 sg13g2_decap_8 FILLER_0_29_194 ();
 sg13g2_decap_8 FILLER_0_29_201 ();
 sg13g2_decap_8 FILLER_0_29_208 ();
 sg13g2_decap_8 FILLER_0_29_215 ();
 sg13g2_decap_8 FILLER_0_29_222 ();
 sg13g2_fill_1 FILLER_0_29_233 ();
 sg13g2_fill_1 FILLER_0_29_249 ();
 sg13g2_decap_8 FILLER_0_30_0 ();
 sg13g2_decap_8 FILLER_0_30_7 ();
 sg13g2_fill_2 FILLER_0_30_14 ();
 sg13g2_fill_1 FILLER_0_30_134 ();
 sg13g2_decap_8 FILLER_0_30_161 ();
 sg13g2_decap_8 FILLER_0_30_168 ();
 sg13g2_decap_8 FILLER_0_30_175 ();
 sg13g2_decap_8 FILLER_0_30_182 ();
 sg13g2_decap_8 FILLER_0_30_189 ();
 sg13g2_decap_8 FILLER_0_30_196 ();
 sg13g2_decap_8 FILLER_0_30_203 ();
 sg13g2_decap_4 FILLER_0_30_210 ();
 sg13g2_fill_1 FILLER_0_30_214 ();
 sg13g2_fill_1 FILLER_0_30_258 ();
 sg13g2_fill_1 FILLER_0_30_267 ();
 sg13g2_fill_1 FILLER_0_30_306 ();
 sg13g2_decap_8 FILLER_0_31_0 ();
 sg13g2_decap_8 FILLER_0_31_7 ();
 sg13g2_decap_8 FILLER_0_31_14 ();
 sg13g2_decap_4 FILLER_0_31_21 ();
 sg13g2_fill_2 FILLER_0_31_25 ();
 sg13g2_fill_2 FILLER_0_31_35 ();
 sg13g2_fill_1 FILLER_0_31_37 ();
 sg13g2_fill_1 FILLER_0_31_76 ();
 sg13g2_fill_2 FILLER_0_31_251 ();
 sg13g2_fill_1 FILLER_0_31_253 ();
 sg13g2_fill_1 FILLER_0_31_258 ();
 sg13g2_fill_2 FILLER_0_31_279 ();
 sg13g2_fill_2 FILLER_0_31_285 ();
 sg13g2_fill_1 FILLER_0_31_293 ();
 sg13g2_fill_1 FILLER_0_31_322 ();
 sg13g2_decap_8 FILLER_0_32_0 ();
 sg13g2_decap_8 FILLER_0_32_7 ();
 sg13g2_decap_8 FILLER_0_32_14 ();
 sg13g2_decap_4 FILLER_0_32_21 ();
 sg13g2_fill_1 FILLER_0_32_25 ();
 sg13g2_fill_1 FILLER_0_32_75 ();
 sg13g2_fill_1 FILLER_0_32_132 ();
 sg13g2_fill_2 FILLER_0_32_138 ();
 sg13g2_fill_2 FILLER_0_32_191 ();
 sg13g2_fill_2 FILLER_0_32_209 ();
 sg13g2_fill_1 FILLER_0_32_211 ();
 sg13g2_fill_2 FILLER_0_32_250 ();
 sg13g2_fill_1 FILLER_0_32_252 ();
 sg13g2_fill_1 FILLER_0_32_307 ();
 sg13g2_fill_1 FILLER_0_32_314 ();
 sg13g2_decap_8 FILLER_0_33_0 ();
 sg13g2_decap_8 FILLER_0_33_7 ();
 sg13g2_decap_8 FILLER_0_33_14 ();
 sg13g2_fill_2 FILLER_0_33_21 ();
 sg13g2_fill_1 FILLER_0_33_23 ();
 sg13g2_fill_2 FILLER_0_33_69 ();
 sg13g2_fill_1 FILLER_0_33_106 ();
 sg13g2_fill_1 FILLER_0_33_142 ();
 sg13g2_fill_1 FILLER_0_33_148 ();
 sg13g2_fill_2 FILLER_0_33_161 ();
 sg13g2_fill_2 FILLER_0_33_279 ();
 sg13g2_fill_1 FILLER_0_33_292 ();
 sg13g2_fill_1 FILLER_0_33_299 ();
 sg13g2_fill_1 FILLER_0_33_309 ();
 sg13g2_decap_8 FILLER_0_34_0 ();
 sg13g2_decap_8 FILLER_0_34_7 ();
 sg13g2_decap_8 FILLER_0_34_14 ();
 sg13g2_decap_4 FILLER_0_34_21 ();
 sg13g2_fill_1 FILLER_0_34_85 ();
 sg13g2_fill_1 FILLER_0_34_90 ();
 sg13g2_fill_1 FILLER_0_34_96 ();
 sg13g2_fill_2 FILLER_0_34_102 ();
 sg13g2_fill_2 FILLER_0_34_109 ();
 sg13g2_fill_2 FILLER_0_34_116 ();
 sg13g2_fill_2 FILLER_0_34_177 ();
 sg13g2_fill_1 FILLER_0_34_183 ();
 sg13g2_fill_1 FILLER_0_34_189 ();
 sg13g2_fill_1 FILLER_0_34_199 ();
 sg13g2_fill_2 FILLER_0_34_228 ();
 sg13g2_fill_1 FILLER_0_34_238 ();
 sg13g2_fill_2 FILLER_0_34_247 ();
 sg13g2_fill_1 FILLER_0_34_253 ();
 sg13g2_fill_2 FILLER_0_34_280 ();
 sg13g2_fill_2 FILLER_0_34_287 ();
 sg13g2_decap_8 FILLER_0_35_0 ();
 sg13g2_decap_8 FILLER_0_35_7 ();
 sg13g2_decap_4 FILLER_0_35_14 ();
 sg13g2_fill_2 FILLER_0_35_18 ();
 sg13g2_fill_1 FILLER_0_35_93 ();
 sg13g2_fill_1 FILLER_0_35_104 ();
 sg13g2_fill_1 FILLER_0_35_136 ();
 sg13g2_fill_2 FILLER_0_35_159 ();
 sg13g2_fill_2 FILLER_0_35_171 ();
 sg13g2_fill_2 FILLER_0_35_204 ();
 sg13g2_fill_1 FILLER_0_35_280 ();
 sg13g2_fill_1 FILLER_0_35_289 ();
 sg13g2_fill_1 FILLER_0_35_295 ();
 sg13g2_fill_2 FILLER_0_35_320 ();
 sg13g2_fill_1 FILLER_0_35_322 ();
 sg13g2_decap_8 FILLER_0_36_0 ();
 sg13g2_decap_8 FILLER_0_36_7 ();
 sg13g2_fill_2 FILLER_0_36_14 ();
 sg13g2_fill_1 FILLER_0_36_16 ();
 sg13g2_fill_2 FILLER_0_36_51 ();
 sg13g2_fill_1 FILLER_0_36_53 ();
 sg13g2_fill_2 FILLER_0_36_68 ();
 sg13g2_fill_1 FILLER_0_36_118 ();
 sg13g2_fill_1 FILLER_0_36_271 ();
 sg13g2_fill_2 FILLER_0_36_294 ();
 sg13g2_fill_1 FILLER_0_36_296 ();
 sg13g2_decap_8 FILLER_0_37_0 ();
 sg13g2_decap_8 FILLER_0_37_7 ();
 sg13g2_decap_4 FILLER_0_37_14 ();
 sg13g2_fill_2 FILLER_0_37_18 ();
 sg13g2_fill_1 FILLER_0_37_66 ();
 sg13g2_fill_1 FILLER_0_37_72 ();
 sg13g2_fill_1 FILLER_0_37_103 ();
 sg13g2_fill_2 FILLER_0_37_108 ();
 sg13g2_fill_1 FILLER_0_37_115 ();
 sg13g2_fill_1 FILLER_0_37_204 ();
 sg13g2_fill_1 FILLER_0_37_238 ();
 sg13g2_decap_8 FILLER_0_38_0 ();
 sg13g2_decap_8 FILLER_0_38_7 ();
 sg13g2_fill_1 FILLER_0_38_14 ();
 sg13g2_decap_4 FILLER_0_38_33 ();
 sg13g2_fill_1 FILLER_0_38_37 ();
 sg13g2_decap_4 FILLER_0_38_45 ();
 sg13g2_fill_1 FILLER_0_38_49 ();
 sg13g2_fill_1 FILLER_0_38_54 ();
 sg13g2_fill_2 FILLER_0_38_108 ();
 sg13g2_fill_1 FILLER_0_38_166 ();
 sg13g2_fill_2 FILLER_0_38_195 ();
 sg13g2_fill_1 FILLER_0_38_230 ();
 sg13g2_fill_2 FILLER_0_38_312 ();
 sg13g2_fill_1 FILLER_0_38_314 ();
 sg13g2_decap_8 FILLER_0_39_0 ();
 sg13g2_decap_8 FILLER_0_39_7 ();
 sg13g2_decap_4 FILLER_0_39_14 ();
 sg13g2_fill_2 FILLER_0_39_114 ();
 sg13g2_fill_1 FILLER_0_39_116 ();
 sg13g2_fill_2 FILLER_0_39_198 ();
 sg13g2_fill_1 FILLER_0_39_288 ();
 sg13g2_fill_1 FILLER_0_39_294 ();
 sg13g2_fill_2 FILLER_0_39_308 ();
 sg13g2_fill_1 FILLER_0_39_310 ();
 sg13g2_decap_8 FILLER_0_40_0 ();
 sg13g2_decap_8 FILLER_0_40_7 ();
 sg13g2_decap_8 FILLER_0_40_14 ();
 sg13g2_decap_4 FILLER_0_40_21 ();
 sg13g2_fill_1 FILLER_0_40_25 ();
 sg13g2_fill_1 FILLER_0_40_81 ();
 sg13g2_fill_1 FILLER_0_40_127 ();
 sg13g2_fill_2 FILLER_0_40_147 ();
 sg13g2_fill_1 FILLER_0_40_153 ();
 sg13g2_fill_2 FILLER_0_40_195 ();
 sg13g2_fill_1 FILLER_0_40_197 ();
 sg13g2_fill_1 FILLER_0_40_288 ();
 sg13g2_fill_2 FILLER_0_40_295 ();
 sg13g2_decap_8 FILLER_0_41_0 ();
 sg13g2_decap_8 FILLER_0_41_7 ();
 sg13g2_decap_8 FILLER_0_41_14 ();
 sg13g2_fill_2 FILLER_0_41_21 ();
 sg13g2_decap_4 FILLER_0_41_40 ();
 sg13g2_fill_2 FILLER_0_41_100 ();
 sg13g2_fill_2 FILLER_0_41_117 ();
 sg13g2_fill_2 FILLER_0_41_159 ();
 sg13g2_fill_1 FILLER_0_41_175 ();
 sg13g2_fill_1 FILLER_0_41_191 ();
 sg13g2_fill_2 FILLER_0_41_208 ();
 sg13g2_fill_1 FILLER_0_41_210 ();
 sg13g2_fill_1 FILLER_0_41_225 ();
 sg13g2_fill_1 FILLER_0_41_236 ();
 sg13g2_fill_2 FILLER_0_41_294 ();
 sg13g2_fill_1 FILLER_0_41_296 ();
 sg13g2_decap_8 FILLER_0_42_0 ();
 sg13g2_decap_8 FILLER_0_42_7 ();
 sg13g2_decap_8 FILLER_0_42_14 ();
 sg13g2_decap_8 FILLER_0_42_21 ();
 sg13g2_decap_8 FILLER_0_42_28 ();
 sg13g2_fill_1 FILLER_0_42_35 ();
 sg13g2_fill_2 FILLER_0_42_73 ();
 sg13g2_fill_2 FILLER_0_42_101 ();
 sg13g2_fill_1 FILLER_0_42_103 ();
 sg13g2_fill_1 FILLER_0_42_143 ();
 sg13g2_fill_2 FILLER_0_42_321 ();
 sg13g2_decap_8 FILLER_0_43_0 ();
 sg13g2_decap_8 FILLER_0_43_7 ();
 sg13g2_decap_8 FILLER_0_43_14 ();
 sg13g2_decap_8 FILLER_0_43_21 ();
 sg13g2_decap_8 FILLER_0_43_28 ();
 sg13g2_decap_4 FILLER_0_43_35 ();
 sg13g2_fill_1 FILLER_0_43_39 ();
 sg13g2_fill_2 FILLER_0_43_129 ();
 sg13g2_fill_2 FILLER_0_43_165 ();
 sg13g2_fill_2 FILLER_0_43_172 ();
 sg13g2_fill_1 FILLER_0_43_174 ();
 sg13g2_fill_2 FILLER_0_43_180 ();
 sg13g2_fill_2 FILLER_0_43_197 ();
 sg13g2_fill_1 FILLER_0_43_208 ();
 sg13g2_fill_2 FILLER_0_43_278 ();
 sg13g2_fill_1 FILLER_0_43_280 ();
 sg13g2_fill_2 FILLER_0_43_291 ();
 sg13g2_fill_1 FILLER_0_43_293 ();
 sg13g2_decap_8 FILLER_0_44_0 ();
 sg13g2_decap_8 FILLER_0_44_7 ();
 sg13g2_decap_8 FILLER_0_44_14 ();
 sg13g2_decap_8 FILLER_0_44_21 ();
 sg13g2_decap_8 FILLER_0_44_28 ();
 sg13g2_decap_4 FILLER_0_44_35 ();
 sg13g2_fill_1 FILLER_0_44_39 ();
 sg13g2_fill_1 FILLER_0_44_112 ();
 sg13g2_fill_1 FILLER_0_44_139 ();
 sg13g2_fill_2 FILLER_0_44_145 ();
 sg13g2_fill_1 FILLER_0_44_152 ();
 sg13g2_fill_2 FILLER_0_44_157 ();
 sg13g2_fill_2 FILLER_0_44_219 ();
 sg13g2_fill_1 FILLER_0_44_221 ();
 sg13g2_fill_1 FILLER_0_44_278 ();
 sg13g2_fill_1 FILLER_0_44_285 ();
 sg13g2_fill_1 FILLER_0_44_299 ();
 sg13g2_fill_2 FILLER_0_44_321 ();
 sg13g2_decap_8 FILLER_0_45_0 ();
 sg13g2_decap_8 FILLER_0_45_7 ();
 sg13g2_decap_8 FILLER_0_45_14 ();
 sg13g2_decap_8 FILLER_0_45_21 ();
 sg13g2_decap_8 FILLER_0_45_28 ();
 sg13g2_decap_4 FILLER_0_45_35 ();
 sg13g2_fill_2 FILLER_0_45_39 ();
 sg13g2_fill_1 FILLER_0_45_77 ();
 sg13g2_fill_2 FILLER_0_45_123 ();
 sg13g2_fill_2 FILLER_0_45_177 ();
 sg13g2_fill_1 FILLER_0_45_185 ();
 sg13g2_fill_1 FILLER_0_45_262 ();
 sg13g2_fill_2 FILLER_0_45_313 ();
 sg13g2_fill_1 FILLER_0_45_315 ();
 sg13g2_decap_8 FILLER_0_46_0 ();
 sg13g2_decap_8 FILLER_0_46_7 ();
 sg13g2_decap_8 FILLER_0_46_14 ();
 sg13g2_decap_8 FILLER_0_46_21 ();
 sg13g2_decap_8 FILLER_0_46_28 ();
 sg13g2_decap_4 FILLER_0_46_35 ();
 sg13g2_fill_1 FILLER_0_46_39 ();
 sg13g2_fill_1 FILLER_0_46_93 ();
 sg13g2_fill_1 FILLER_0_46_147 ();
 sg13g2_fill_1 FILLER_0_46_153 ();
 sg13g2_fill_1 FILLER_0_46_180 ();
 sg13g2_fill_1 FILLER_0_46_186 ();
 sg13g2_fill_2 FILLER_0_46_230 ();
 sg13g2_fill_1 FILLER_0_46_268 ();
 sg13g2_fill_2 FILLER_0_46_315 ();
 sg13g2_fill_1 FILLER_0_46_317 ();
 sg13g2_decap_8 FILLER_0_47_0 ();
 sg13g2_fill_2 FILLER_0_47_7 ();
 sg13g2_fill_1 FILLER_0_47_47 ();
 sg13g2_decap_4 FILLER_0_47_64 ();
 sg13g2_fill_2 FILLER_0_47_104 ();
 sg13g2_fill_2 FILLER_0_47_114 ();
 sg13g2_fill_1 FILLER_0_47_175 ();
 sg13g2_fill_1 FILLER_0_47_223 ();
 sg13g2_fill_1 FILLER_0_47_256 ();
 sg13g2_fill_1 FILLER_0_47_263 ();
 sg13g2_fill_2 FILLER_0_47_269 ();
 sg13g2_fill_1 FILLER_0_47_271 ();
 sg13g2_fill_1 FILLER_0_47_296 ();
 sg13g2_fill_1 FILLER_0_47_312 ();
 sg13g2_fill_2 FILLER_0_47_320 ();
 sg13g2_fill_1 FILLER_0_47_322 ();
 sg13g2_decap_8 FILLER_0_48_0 ();
 sg13g2_decap_8 FILLER_0_48_7 ();
 sg13g2_fill_2 FILLER_0_48_14 ();
 sg13g2_fill_1 FILLER_0_48_16 ();
 sg13g2_decap_8 FILLER_0_48_21 ();
 sg13g2_decap_8 FILLER_0_48_28 ();
 sg13g2_decap_8 FILLER_0_48_35 ();
 sg13g2_decap_8 FILLER_0_48_42 ();
 sg13g2_fill_1 FILLER_0_48_49 ();
 sg13g2_fill_2 FILLER_0_48_71 ();
 sg13g2_fill_2 FILLER_0_48_100 ();
 sg13g2_fill_1 FILLER_0_48_102 ();
 sg13g2_fill_1 FILLER_0_48_137 ();
 sg13g2_fill_2 FILLER_0_48_193 ();
 sg13g2_fill_1 FILLER_0_48_268 ();
 sg13g2_fill_1 FILLER_0_48_273 ();
 sg13g2_decap_8 FILLER_0_49_0 ();
 sg13g2_decap_8 FILLER_0_49_7 ();
 sg13g2_decap_8 FILLER_0_49_14 ();
 sg13g2_decap_8 FILLER_0_49_21 ();
 sg13g2_decap_8 FILLER_0_49_28 ();
 sg13g2_fill_1 FILLER_0_49_35 ();
 sg13g2_fill_2 FILLER_0_49_105 ();
 sg13g2_fill_1 FILLER_0_49_145 ();
 sg13g2_fill_1 FILLER_0_49_179 ();
 sg13g2_fill_2 FILLER_0_49_203 ();
 sg13g2_fill_1 FILLER_0_49_205 ();
 sg13g2_fill_1 FILLER_0_49_221 ();
 sg13g2_fill_2 FILLER_0_49_231 ();
 sg13g2_decap_8 FILLER_0_50_0 ();
 sg13g2_decap_8 FILLER_0_50_7 ();
 sg13g2_decap_8 FILLER_0_50_14 ();
 sg13g2_decap_8 FILLER_0_50_21 ();
 sg13g2_fill_2 FILLER_0_50_28 ();
 sg13g2_fill_1 FILLER_0_50_65 ();
 sg13g2_fill_1 FILLER_0_50_96 ();
 sg13g2_fill_2 FILLER_0_50_106 ();
 sg13g2_fill_1 FILLER_0_50_150 ();
 sg13g2_fill_1 FILLER_0_50_215 ();
 sg13g2_fill_1 FILLER_0_50_296 ();
 sg13g2_decap_8 FILLER_0_51_0 ();
 sg13g2_decap_8 FILLER_0_51_7 ();
 sg13g2_decap_8 FILLER_0_51_14 ();
 sg13g2_decap_8 FILLER_0_51_21 ();
 sg13g2_decap_8 FILLER_0_51_28 ();
 sg13g2_fill_1 FILLER_0_51_35 ();
 sg13g2_fill_2 FILLER_0_51_116 ();
 sg13g2_fill_1 FILLER_0_51_156 ();
 sg13g2_fill_1 FILLER_0_51_171 ();
 sg13g2_fill_2 FILLER_0_51_282 ();
 sg13g2_fill_1 FILLER_0_51_306 ();
 sg13g2_fill_2 FILLER_0_51_321 ();
 sg13g2_decap_8 FILLER_0_52_4 ();
 sg13g2_decap_8 FILLER_0_52_11 ();
 sg13g2_decap_8 FILLER_0_52_18 ();
 sg13g2_fill_1 FILLER_0_52_25 ();
 sg13g2_fill_2 FILLER_0_52_169 ();
 sg13g2_fill_2 FILLER_0_52_201 ();
 sg13g2_fill_2 FILLER_0_52_253 ();
 sg13g2_fill_1 FILLER_0_52_298 ();
 sg13g2_fill_2 FILLER_0_52_309 ();
 sg13g2_fill_2 FILLER_0_52_321 ();
 sg13g2_fill_2 FILLER_0_53_0 ();
 sg13g2_fill_1 FILLER_0_53_2 ();
 sg13g2_fill_1 FILLER_0_53_7 ();
 sg13g2_decap_4 FILLER_0_53_16 ();
 sg13g2_fill_1 FILLER_0_53_20 ();
 sg13g2_fill_1 FILLER_0_53_75 ();
 sg13g2_fill_2 FILLER_0_53_80 ();
 sg13g2_fill_2 FILLER_0_53_155 ();
 sg13g2_fill_1 FILLER_0_53_205 ();
 sg13g2_fill_2 FILLER_0_53_215 ();
 sg13g2_fill_1 FILLER_0_54_0 ();
 sg13g2_fill_1 FILLER_0_54_28 ();
 sg13g2_fill_1 FILLER_0_54_82 ();
 sg13g2_fill_1 FILLER_0_54_103 ();
 sg13g2_fill_2 FILLER_0_54_120 ();
 sg13g2_fill_1 FILLER_0_54_122 ();
 sg13g2_fill_1 FILLER_0_54_127 ();
 sg13g2_fill_1 FILLER_0_54_132 ();
 sg13g2_fill_1 FILLER_0_54_141 ();
 sg13g2_fill_1 FILLER_0_54_167 ();
 sg13g2_fill_1 FILLER_0_54_250 ();
 sg13g2_fill_2 FILLER_0_54_279 ();
 sg13g2_fill_1 FILLER_0_54_281 ();
 sg13g2_fill_1 FILLER_0_54_287 ();
 sg13g2_fill_1 FILLER_0_54_306 ();
 sg13g2_fill_2 FILLER_0_54_321 ();
 sg13g2_fill_2 FILLER_0_55_40 ();
 sg13g2_fill_1 FILLER_0_55_161 ();
 sg13g2_fill_2 FILLER_0_55_188 ();
 sg13g2_fill_1 FILLER_0_55_199 ();
 sg13g2_fill_2 FILLER_0_55_253 ();
 sg13g2_fill_2 FILLER_0_55_315 ();
 sg13g2_fill_1 FILLER_0_55_322 ();
 sg13g2_fill_2 FILLER_0_56_4 ();
 sg13g2_fill_1 FILLER_0_56_6 ();
 sg13g2_fill_1 FILLER_0_56_75 ();
 sg13g2_fill_2 FILLER_0_56_293 ();
 sg13g2_fill_2 FILLER_0_56_321 ();
 sg13g2_fill_2 FILLER_0_57_76 ();
 sg13g2_fill_2 FILLER_0_57_154 ();
 sg13g2_fill_1 FILLER_0_57_160 ();
 sg13g2_fill_1 FILLER_0_57_166 ();
 sg13g2_fill_1 FILLER_0_57_171 ();
 sg13g2_fill_1 FILLER_0_57_176 ();
 sg13g2_fill_2 FILLER_0_57_211 ();
 sg13g2_fill_2 FILLER_0_57_217 ();
 sg13g2_fill_1 FILLER_0_57_318 ();
 assign uio_oe[0] = net101;
 assign uio_oe[7] = net98;
endmodule
